module test_07 (N1, N2, N3, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39);

input N1; 
input N2; 
input N3; 

output N26; 
output N27; 
output N28; 
output N29; 
output N30; 
output N31; 
output N32; 
output N33; 
output N34; 
output N35; 
output N36; 
output N37; 
output N38; 
output N39; 

wire N4; 
wire N5; 
wire N6; 
wire N7; 
wire N8; 
wire N9; 
wire N10; 
wire N11; 
wire N12; 
wire N13; 
wire N14; 
wire N15; 
wire N16; 
wire N17; 
wire N18; 
wire N19; 
wire N20; 
wire N21; 
wire N22; 
wire N23; 
wire N24; 
wire N25; 

assign N4 = ~(N2); 
assign N5 = ~(N3); 
assign N6 = N2 & N1; 
assign N7 = ~(N2); 
assign N8 = ~(N2); 
assign N9 = ~(N1); 
assign N10 = ~(N5); 
assign N11 = ~(N6); 
assign N12 = ~(N2); 
assign N13 = N4 | N9; 
assign N14 = N9 | N3; 
assign N15 = ~(N3); 
assign N16 = N6 | N9 | N8 | N1 | N3 | N5 | N2 | N7 | N4; 
assign N17 = ~(N9); 
assign N18 = N3 | N9; 
assign N19 = N16 & N4; 
assign N20 = N8 | N4; 
assign N21 = N12 & N17; 
assign N22 = ~(N19); 
assign N23 = N1 & N13 & N6; 
assign N24 = N7 & N19 & N20 & N8; 
assign N25 = N15 | N7; 
assign N26 = ~(N21); 
assign N27 = N6 & N18 & N23; 
assign N28 = ~(N22); 
assign N29 = N4 & N19 & N10 & N16 & N3 & N11 & N6 & N17 & N23; 
assign N30 = ~(N11); 
assign N31 = ~(N10); 
assign N32 = ~(N14); 
assign N33 = N19 | N24 | N16 | N11 | N13 | N5 | N25 | N1 | N8; 
assign N34 = N19 & N9 & N22 & N21 & N18 & N20 & N24 & N25 & N1; 
assign N35 = ~(N5); 
assign N36 = ~(N25); 
assign N37 = N21 | N20 | N7 | N13 | N22 | N11 | N16 | N23 | N5; 
assign N38 = N11 | N21 | N13 | N4 | N24 | N20 | N18 | N5 | N25; 
assign N39 = ~(N24); 
endmodule
