module test_03 (N1, N2, N3, N4, N5, N32, N33, N34, N35, N36, N37, N38);

input N1; 
input N2; 
input N3; 
input N4; 
input N5; 

output N32; 
output N33; 
output N34; 
output N35; 
output N36; 
output N37; 
output N38; 

wire N6; 
wire N7; 
wire N8; 
wire N9; 
wire N10; 
wire N11; 
wire N12; 
wire N13; 
wire N14; 
wire N15; 
wire N16; 
wire N17; 
wire N18; 
wire N19; 
wire N20; 
wire N21; 
wire N22; 
wire N23; 
wire N24; 
wire N25; 
wire N26; 
wire N27; 
wire N28; 
wire N29; 
wire N30; 
wire N31; 

assign N6 = ~(N4); 
assign N7 = ~(N3); 
assign N8 = ~(N1); 
assign N9 = ~(N3); 
assign N10 = ~(N1); 
assign N11 = ~(N2); 
assign N12 = ~(N7); 
assign N13 = ~(N3); 
assign N14 = N1 | N8 | N10; 
assign N15 = ~(N10); 
assign N16 = N7 & N9; 
assign N17 = ~(N2); 
assign N18 = N14 & N12; 
assign N19 = N6 | N10; 
assign N20 = ~(N16); 
assign N21 = N12 & N8; 
assign N22 = ~(N10); 
assign N23 = N18 | N20 | N17; 
assign N24 = N15 & N12; 
assign N25 = N5 & N17 & N19 & N15; 
assign N26 = ~(N6); 
assign N27 = ~(N21); 
assign N28 = N4 | N16 | N22 | N2; 
assign N29 = ~(N26); 
assign N30 = ~(N5); 
assign N31 = N21 & N25 & N6; 
assign N32 = ~(N31); 
assign N33 = N2 | N28 | N30; 
assign N34 = N18 | N16 | N26 | N23 | N28 | N14 | N5 | N24 | N9; 
assign N35 = N11 | N13; 
assign N36 = N24 | N29; 
assign N37 = N10 & N23; 
assign N38 = N9 | N27; 
endmodule
