module test_09 (N1, N2, N3, N4, N5, N6, N7, N32, N33, N34, N35, N36, N37, N38);

input N1; 
input N2; 
input N3; 
input N4; 
input N5; 
input N6; 
input N7; 

output N32; 
output N33; 
output N34; 
output N35; 
output N36; 
output N37; 
output N38; 

wire N8; 
wire N9; 
wire N10; 
wire N11; 
wire N12; 
wire N13; 
wire N14; 
wire N15; 
wire N16; 
wire N17; 
wire N18; 
wire N19; 
wire N20; 
wire N21; 
wire N22; 
wire N23; 
wire N24; 
wire N25; 
wire N26; 
wire N27; 
wire N28; 
wire N29; 
wire N30; 
wire N31; 

assign N8 = ~(N1); 
assign N9 = N5 & N4; 
assign N10 = N4 & N2; 
assign N11 = ~(N4); 
assign N12 = ~(N9); 
assign N13 = N2 | N1; 
assign N14 = ~(N12); 
assign N15 = ~(N10); 
assign N16 = N6 & N11; 
assign N17 = ~(N16); 
assign N18 = ~(N9); 
assign N19 = N9 | N11; 
assign N20 = N7 & N14 & N15; 
assign N21 = ~(N1); 
assign N22 = N16 & N5; 
assign N23 = N1 & N17 & N14; 
assign N24 = ~(N10); 
assign N25 = N8 | N10 | N11 | N20 | N22; 
assign N26 = N13 & N21; 
assign N27 = ~(N16); 
assign N28 = N23 & N27; 
assign N29 = N21 & N13; 
assign N30 = ~(N10); 
assign N31 = N3 | N15 | N25; 
assign N32 = ~(N31); 
assign N33 = ~(N29); 
assign N34 = N19 | N30; 
assign N35 = N24 | N28; 
assign N36 = N18 & N25; 
assign N37 = ~(N27); 
assign N38 = ~(N26); 
endmodule
