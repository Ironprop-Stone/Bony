module Depth_10_20_Nodes_200_400_S002 (N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341, N342, N343, N344);

input N1; 
input N2; 
input N3; 
input N4; 
input N5; 
input N6; 
input N7; 
input N8; 
input N9; 
input N10; 

output N331; 
output N332; 
output N333; 
output N334; 
output N335; 
output N336; 
output N337; 
output N338; 
output N339; 
output N340; 
output N341; 
output N342; 
output N343; 
output N344; 

wire N11; 
wire N12; 
wire N13; 
wire N14; 
wire N15; 
wire N16; 
wire N17; 
wire N18; 
wire N19; 
wire N20; 
wire N21; 
wire N22; 
wire N23; 
wire N24; 
wire N25; 
wire N26; 
wire N27; 
wire N28; 
wire N29; 
wire N30; 
wire N31; 
wire N32; 
wire N33; 
wire N34; 
wire N35; 
wire N36; 
wire N37; 
wire N38; 
wire N39; 
wire N40; 
wire N41; 
wire N42; 
wire N43; 
wire N44; 
wire N45; 
wire N46; 
wire N47; 
wire N48; 
wire N49; 
wire N50; 
wire N51; 
wire N52; 
wire N53; 
wire N54; 
wire N55; 
wire N56; 
wire N57; 
wire N58; 
wire N59; 
wire N60; 
wire N61; 
wire N62; 
wire N63; 
wire N64; 
wire N65; 
wire N66; 
wire N67; 
wire N68; 
wire N69; 
wire N70; 
wire N71; 
wire N72; 
wire N73; 
wire N74; 
wire N75; 
wire N76; 
wire N77; 
wire N78; 
wire N79; 
wire N80; 
wire N81; 
wire N82; 
wire N83; 
wire N84; 
wire N85; 
wire N86; 
wire N87; 
wire N88; 
wire N89; 
wire N90; 
wire N91; 
wire N92; 
wire N93; 
wire N94; 
wire N95; 
wire N96; 
wire N97; 
wire N98; 
wire N99; 
wire N100; 
wire N101; 
wire N102; 
wire N103; 
wire N104; 
wire N105; 
wire N106; 
wire N107; 
wire N108; 
wire N109; 
wire N110; 
wire N111; 
wire N112; 
wire N113; 
wire N114; 
wire N115; 
wire N116; 
wire N117; 
wire N118; 
wire N119; 
wire N120; 
wire N121; 
wire N122; 
wire N123; 
wire N124; 
wire N125; 
wire N126; 
wire N127; 
wire N128; 
wire N129; 
wire N130; 
wire N131; 
wire N132; 
wire N133; 
wire N134; 
wire N135; 
wire N136; 
wire N137; 
wire N138; 
wire N139; 
wire N140; 
wire N141; 
wire N142; 
wire N143; 
wire N144; 
wire N145; 
wire N146; 
wire N147; 
wire N148; 
wire N149; 
wire N150; 
wire N151; 
wire N152; 
wire N153; 
wire N154; 
wire N155; 
wire N156; 
wire N157; 
wire N158; 
wire N159; 
wire N160; 
wire N161; 
wire N162; 
wire N163; 
wire N164; 
wire N165; 
wire N166; 
wire N167; 
wire N168; 
wire N169; 
wire N170; 
wire N171; 
wire N172; 
wire N173; 
wire N174; 
wire N175; 
wire N176; 
wire N177; 
wire N178; 
wire N179; 
wire N180; 
wire N181; 
wire N182; 
wire N183; 
wire N184; 
wire N185; 
wire N186; 
wire N187; 
wire N188; 
wire N189; 
wire N190; 
wire N191; 
wire N192; 
wire N193; 
wire N194; 
wire N195; 
wire N196; 
wire N197; 
wire N198; 
wire N199; 
wire N200; 
wire N201; 
wire N202; 
wire N203; 
wire N204; 
wire N205; 
wire N206; 
wire N207; 
wire N208; 
wire N209; 
wire N210; 
wire N211; 
wire N212; 
wire N213; 
wire N214; 
wire N215; 
wire N216; 
wire N217; 
wire N218; 
wire N219; 
wire N220; 
wire N221; 
wire N222; 
wire N223; 
wire N224; 
wire N225; 
wire N226; 
wire N227; 
wire N228; 
wire N229; 
wire N230; 
wire N231; 
wire N232; 
wire N233; 
wire N234; 
wire N235; 
wire N236; 
wire N237; 
wire N238; 
wire N239; 
wire N240; 
wire N241; 
wire N242; 
wire N243; 
wire N244; 
wire N245; 
wire N246; 
wire N247; 
wire N248; 
wire N249; 
wire N250; 
wire N251; 
wire N252; 
wire N253; 
wire N254; 
wire N255; 
wire N256; 
wire N257; 
wire N258; 
wire N259; 
wire N260; 
wire N261; 
wire N262; 
wire N263; 
wire N264; 
wire N265; 
wire N266; 
wire N267; 
wire N268; 
wire N269; 
wire N270; 
wire N271; 
wire N272; 
wire N273; 
wire N274; 
wire N275; 
wire N276; 
wire N277; 
wire N278; 
wire N279; 
wire N280; 
wire N281; 
wire N282; 
wire N283; 
wire N284; 
wire N285; 
wire N286; 
wire N287; 
wire N288; 
wire N289; 
wire N290; 
wire N291; 
wire N292; 
wire N293; 
wire N294; 
wire N295; 
wire N296; 
wire N297; 
wire N298; 
wire N299; 
wire N300; 
wire N301; 
wire N302; 
wire N303; 
wire N304; 
wire N305; 
wire N306; 
wire N307; 
wire N308; 
wire N309; 
wire N310; 
wire N311; 
wire N312; 
wire N313; 
wire N314; 
wire N315; 
wire N316; 
wire N317; 
wire N318; 
wire N319; 
wire N320; 
wire N321; 
wire N322; 
wire N323; 
wire N324; 
wire N325; 
wire N326; 
wire N327; 
wire N328; 
wire N329; 
wire N330; 

assign N11 = ~(N4); 
assign N12 = ~(N3); 
assign N13 = ~(N2); 
assign N14 = ~(N8); 
assign N15 = ~(N2); 
assign N16 = ~(N4); 
assign N17 = ~(N10); 
assign N18 = ~(N8); 
assign N19 = ~(N8); 
assign N20 = ~(N3); 
assign N21 = N6 | N9 | N5; 
assign N22 = ~(N2); 
assign N23 = ~(N19); 
assign N24 = ~(N21); 
assign N25 = ~(N5); 
assign N26 = ~(N22); 
assign N27 = ~(N8); 
assign N28 = N15 & N4; 
assign N29 = ~(N22); 
assign N30 = ~(N16); 
assign N31 = ~(N14); 
assign N32 = ~(N7); 
assign N33 = ~(N14); 
assign N34 = ~(N16); 
assign N35 = ~(N21); 
assign N36 = N32 & N12; 
assign N37 = N5 | N17; 
assign N38 = ~(N18); 
assign N39 = ~(N34); 
assign N40 = ~(N21); 
assign N41 = ~(N11); 
assign N42 = ~(N7); 
assign N43 = ~(N26); 
assign N44 = ~(N2); 
assign N45 = ~(N36); 
assign N46 = ~(N7); 
assign N47 = N30 | N12; 
assign N48 = N2 | N29; 
assign N49 = N22 & N30; 
assign N50 = N16 & N41; 
assign N51 = N7 | N28 | N22; 
assign N52 = ~(N6); 
assign N53 = ~(N4); 
assign N54 = ~(N5); 
assign N55 = ~(N40); 
assign N56 = N14 | N47; 
assign N57 = ~(N31); 
assign N58 = N43 | N32; 
assign N59 = ~(N34); 
assign N60 = ~(N47); 
assign N61 = ~(N26); 
assign N62 = ~(N26); 
assign N63 = N52 & N40; 
assign N64 = N3 | N27; 
assign N65 = ~(N19); 
assign N66 = N49 & N48; 
assign N67 = N47 & N29; 
assign N68 = ~(N37); 
assign N69 = N25 | N41; 
assign N70 = N40 & N9; 
assign N71 = ~(N41); 
assign N72 = ~(N35); 
assign N73 = ~(N40); 
assign N74 = N27 | N31; 
assign N75 = ~(N36); 
assign N76 = ~(N38); 
assign N77 = ~(N38); 
assign N78 = ~(N39); 
assign N79 = ~(N15); 
assign N80 = ~(N3); 
assign N81 = N10 | N37; 
assign N82 = ~(N28); 
assign N83 = ~(N73); 
assign N84 = ~(N37); 
assign N85 = ~(N49); 
assign N86 = ~(N49); 
assign N87 = N70 | N19; 
assign N88 = ~(N55); 
assign N89 = ~(N18); 
assign N90 = ~(N36); 
assign N91 = N36 | N24; 
assign N92 = ~(N44); 
assign N93 = ~(N39); 
assign N94 = ~(N14); 
assign N95 = N54 & N20; 
assign N96 = ~(N38); 
assign N97 = ~(N36); 
assign N98 = ~(N54); 
assign N99 = N17 | N21; 
assign N100 = ~(N35); 
assign N101 = ~(N55); 
assign N102 = ~(N43); 
assign N103 = ~(N6); 
assign N104 = ~(N15); 
assign N105 = ~(N47); 
assign N106 = ~(N22); 
assign N107 = ~(N14); 
assign N108 = ~(N50); 
assign N109 = ~(N59); 
assign N110 = ~(N5); 
assign N111 = ~(N61); 
assign N112 = ~(N41); 
assign N113 = ~(N6); 
assign N114 = ~(N6); 
assign N115 = ~(N40); 
assign N116 = ~(N43); 
assign N117 = ~(N72); 
assign N118 = ~(N42); 
assign N119 = ~(N13); 
assign N120 = ~(N34); 
assign N121 = ~(N36); 
assign N122 = ~(N73); 
assign N123 = ~(N17); 
assign N124 = N8 & N99 & N68; 
assign N125 = ~(N58); 
assign N126 = N46 | N19; 
assign N127 = N80 | N20; 
assign N128 = N63 | N15; 
assign N129 = N26 | N60 | N77 | N7; 
assign N130 = N71 & N15; 
assign N131 = N68 & N90 & N101 & N70; 
assign N132 = ~(N29); 
assign N133 = N58 | N84 | N49; 
assign N134 = N18 & N29 & N69; 
assign N135 = ~(N72); 
assign N136 = N21 & N26; 
assign N137 = N51 | N83 | N53; 
assign N138 = ~(N46); 
assign N139 = N31 | N88 | N71; 
assign N140 = N39 | N70; 
assign N141 = ~(N86); 
assign N142 = ~(N13); 
assign N143 = N1 | N12 | N134; 
assign N144 = ~(N13); 
assign N145 = ~(N131); 
assign N146 = ~(N34); 
assign N147 = ~(N132); 
assign N148 = ~(N133); 
assign N149 = ~(N28); 
assign N150 = N129 & N10; 
assign N151 = ~(N39); 
assign N152 = N73 & N109 & N62; 
assign N153 = N4 & N33 & N43; 
assign N154 = ~(N132); 
assign N155 = ~(N28); 
assign N156 = N50 | N125 | N131 | N66; 
assign N157 = N119 & N129; 
assign N158 = ~(N97); 
assign N159 = ~(N55); 
assign N160 = N137 & N29; 
assign N161 = ~(N50); 
assign N162 = ~(N17); 
assign N163 = ~(N32); 
assign N164 = N44 | N46; 
assign N165 = ~(N3); 
assign N166 = ~(N59); 
assign N167 = N56 & N66 & N59; 
assign N168 = N24 | N160 | N162; 
assign N169 = N45 & N150; 
assign N170 = N42 & N141; 
assign N171 = N35 & N78 & N114 & N132 & N137; 
assign N172 = N19 & N107 & N118; 
assign N173 = ~(N23); 
assign N174 = N11 | N13 | N20 | N61 | N86 | N108 | N41; 
assign N175 = ~(N51); 
assign N176 = ~(N16); 
assign N177 = ~(N27); 
assign N178 = ~(N20); 
assign N179 = ~(N128); 
assign N180 = ~(N13); 
assign N181 = ~(N128); 
assign N182 = N75 | N38; 
assign N183 = ~(N17); 
assign N184 = N100 | N172 | N138; 
assign N185 = ~(N43); 
assign N186 = ~(N33); 
assign N187 = ~(N137); 
assign N188 = ~(N42); 
assign N189 = ~(N34); 
assign N190 = N140 | N20; 
assign N191 = ~(N161); 
assign N192 = N62 & N72 & N58; 
assign N193 = ~(N17); 
assign N194 = N37 | N79 | N65; 
assign N195 = ~(N168); 
assign N196 = N69 & N132; 
assign N197 = ~(N25); 
assign N198 = N142 & N61; 
assign N199 = ~(N30); 
assign N200 = N113 & N52; 
assign N201 = ~(N128); 
assign N202 = N166 | N93; 
assign N203 = ~(N28); 
assign N204 = N41 | N35; 
assign N205 = ~(N38); 
assign N206 = N85 & N128 & N135; 
assign N207 = ~(N72); 
assign N208 = N57 | N97; 
assign N209 = ~(N60); 
assign N210 = ~(N102); 
assign N211 = ~(N4); 
assign N212 = ~(N209); 
assign N213 = ~(N101); 
assign N214 = N38 & N48 & N53 & N182 & N198 & N98; 
assign N215 = N105 | N47; 
assign N216 = N55 | N92 | N117 | N133 | N78; 
assign N217 = N179 | N7; 
assign N218 = N115 & N72; 
assign N219 = N110 & N95; 
assign N220 = N201 & N23; 
assign N221 = N196 & N102; 
assign N222 = N93 & N103; 
assign N223 = N136 & N164 & N80; 
assign N224 = ~(N74); 
assign N225 = ~(N116); 
assign N226 = ~(N10); 
assign N227 = ~(N157); 
assign N228 = ~(N23); 
assign N229 = N96 & N115; 
assign N230 = ~(N66); 
assign N231 = ~(N33); 
assign N232 = N103 & N192 & N37; 
assign N233 = ~(N50); 
assign N234 = N120 & N144 & N202 & N18; 
assign N235 = ~(N147); 
assign N236 = ~(N60); 
assign N237 = ~(N71); 
assign N238 = N127 | N139; 
assign N239 = ~(N207); 
assign N240 = N67 & N73; 
assign N241 = ~(N188); 
assign N242 = ~(N108); 
assign N243 = N112 | N87; 
assign N244 = N183 & N18; 
assign N245 = ~(N39); 
assign N246 = ~(N72); 
assign N247 = ~(N39); 
assign N248 = ~(N112); 
assign N249 = ~(N15); 
assign N250 = N190 | N86; 
assign N251 = ~(N130); 
assign N252 = ~(N129); 
assign N253 = N163 | N219 | N134; 
assign N254 = ~(N128); 
assign N255 = ~(N65); 
assign N256 = N76 & N60; 
assign N257 = N116 & N33; 
assign N258 = ~(N171); 
assign N259 = N173 & N35; 
assign N260 = N89 & N131; 
assign N261 = N139 & N81; 
assign N262 = N65 | N130 | N199 | N105; 
assign N263 = N98 | N102 | N123 | N185 | N222 | N224; 
assign N264 = N64 | N135 | N143 | N161 | N194 | N95; 
assign N265 = N82 & N147 & N229 & N251 & N32; 
assign N266 = N91 & N126 & N152 & N189 & N240 & N30; 
assign N267 = N111 | N124 | N134 | N215 | N10; 
assign N268 = N148 | N211 | N131; 
assign N269 = N106 & N149 & N153 & N235 & N98; 
assign N270 = N175 | N264 | N136; 
assign N271 = N230 | N245 | N70; 
assign N272 = ~(N99); 
assign N273 = N81 | N95 | N97 | N169 | N177 | N243 | N263 | N52; 
assign N274 = N94 | N121 | N195 | N231 | N137; 
assign N275 = N228 | N237 | N244; 
assign N276 = N87 & N138 & N239 & N265 & N119; 
assign N277 = N104 | N217 | N69; 
assign N278 = ~(N16); 
assign N279 = ~(N104); 
assign N280 = N167 & N59; 
assign N281 = ~(N79); 
assign N282 = N187 | N276 | N125; 
assign N283 = ~(N27); 
assign N284 = N157 & N22; 
assign N285 = ~(N147); 
assign N286 = ~(N221); 
assign N287 = N180 & N250; 
assign N288 = N170 & N11; 
assign N289 = N221 | N247 | N1; 
assign N290 = N176 & N1; 
assign N291 = ~(N75); 
assign N292 = N145 | N273; 
assign N293 = N216 & N254 & N28; 
assign N294 = ~(N49); 
assign N295 = ~(N122); 
assign N296 = ~(N203); 
assign N297 = N156 | N269; 
assign N298 = ~(N108); 
assign N299 = N151 & N234 & N246 & N267 & N9; 
assign N300 = N258 & N66; 
assign N301 = N283 | N43; 
assign N302 = N186 | N293 | N100; 
assign N303 = N226 | N242 | N270 | N279 | N141; 
assign N304 = N174 | N212 | N255; 
assign N305 = N277 | N94; 
assign N306 = N214 | N252 | N268 | N298 | N25; 
assign N307 = ~(N158); 
assign N308 = ~(N287); 
assign N309 = N146 | N165 | N233 | N241 | N249 | N253; 
assign N310 = ~(N213); 
assign N311 = N218 | N232 | N286; 
assign N312 = N154 & N291 & N92; 
assign N313 = N159 | N129; 
assign N314 = N184 | N271; 
assign N315 = N168 & N191 & N223 & N287 & N46; 
assign N316 = N155 | N200 | N85; 
assign N317 = ~(N135); 
assign N318 = ~(N61); 
assign N319 = ~(N225); 
assign N320 = N257 & N262 & N275 & N46; 
assign N321 = N197 & N205; 
assign N322 = ~(N296); 
assign N323 = ~(N207); 
assign N324 = N238 & N259 & N260 & N302; 
assign N325 = N288 & N290 & N98; 
assign N326 = N210 & N313 & N141; 
assign N327 = N206 | N220 | N316; 
assign N328 = N181 & N208 & N304 & N309; 
assign N329 = N284 | N11; 
assign N330 = N193 & N272 & N294; 
assign N331 = N281 | N289 | N318; 
assign N332 = N261 & N328; 
assign N333 = N278 & N299 & N306 & N322 & N325; 
assign N334 = N319 | N323 | N326 | N327 | N329; 
assign N335 = N292 & N320; 
assign N336 = ~(N305); 
assign N337 = N282 | N308; 
assign N338 = N225 | N280 | N297 | N303 | N310 | N321; 
assign N339 = N178 & N295 & N330; 
assign N340 = N204 | N248 | N285 | N314 | N324; 
assign N341 = N256 & N266 & N274 & N312; 
assign N342 = ~(N311); 
assign N343 = N236 & N301 & N307 & N315; 
assign N344 = N227 | N300 | N317; 
endmodule
