module Depth_10_20_Nodes_200_400_S006 (N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N445, N446, N447, N448, N449, N450, N451, N452, N453, N454, N455, N456, N457, N458, N459, N460, N461, N462, N463, N464, N465, N466, N467, N468, N469, N470, N471);

input N1; 
input N2; 
input N3; 
input N4; 
input N5; 
input N6; 
input N7; 
input N8; 
input N9; 
input N10; 
input N11; 
input N12; 
input N13; 

output N445; 
output N446; 
output N447; 
output N448; 
output N449; 
output N450; 
output N451; 
output N452; 
output N453; 
output N454; 
output N455; 
output N456; 
output N457; 
output N458; 
output N459; 
output N460; 
output N461; 
output N462; 
output N463; 
output N464; 
output N465; 
output N466; 
output N467; 
output N468; 
output N469; 
output N470; 
output N471; 

wire N14; 
wire N15; 
wire N16; 
wire N17; 
wire N18; 
wire N19; 
wire N20; 
wire N21; 
wire N22; 
wire N23; 
wire N24; 
wire N25; 
wire N26; 
wire N27; 
wire N28; 
wire N29; 
wire N30; 
wire N31; 
wire N32; 
wire N33; 
wire N34; 
wire N35; 
wire N36; 
wire N37; 
wire N38; 
wire N39; 
wire N40; 
wire N41; 
wire N42; 
wire N43; 
wire N44; 
wire N45; 
wire N46; 
wire N47; 
wire N48; 
wire N49; 
wire N50; 
wire N51; 
wire N52; 
wire N53; 
wire N54; 
wire N55; 
wire N56; 
wire N57; 
wire N58; 
wire N59; 
wire N60; 
wire N61; 
wire N62; 
wire N63; 
wire N64; 
wire N65; 
wire N66; 
wire N67; 
wire N68; 
wire N69; 
wire N70; 
wire N71; 
wire N72; 
wire N73; 
wire N74; 
wire N75; 
wire N76; 
wire N77; 
wire N78; 
wire N79; 
wire N80; 
wire N81; 
wire N82; 
wire N83; 
wire N84; 
wire N85; 
wire N86; 
wire N87; 
wire N88; 
wire N89; 
wire N90; 
wire N91; 
wire N92; 
wire N93; 
wire N94; 
wire N95; 
wire N96; 
wire N97; 
wire N98; 
wire N99; 
wire N100; 
wire N101; 
wire N102; 
wire N103; 
wire N104; 
wire N105; 
wire N106; 
wire N107; 
wire N108; 
wire N109; 
wire N110; 
wire N111; 
wire N112; 
wire N113; 
wire N114; 
wire N115; 
wire N116; 
wire N117; 
wire N118; 
wire N119; 
wire N120; 
wire N121; 
wire N122; 
wire N123; 
wire N124; 
wire N125; 
wire N126; 
wire N127; 
wire N128; 
wire N129; 
wire N130; 
wire N131; 
wire N132; 
wire N133; 
wire N134; 
wire N135; 
wire N136; 
wire N137; 
wire N138; 
wire N139; 
wire N140; 
wire N141; 
wire N142; 
wire N143; 
wire N144; 
wire N145; 
wire N146; 
wire N147; 
wire N148; 
wire N149; 
wire N150; 
wire N151; 
wire N152; 
wire N153; 
wire N154; 
wire N155; 
wire N156; 
wire N157; 
wire N158; 
wire N159; 
wire N160; 
wire N161; 
wire N162; 
wire N163; 
wire N164; 
wire N165; 
wire N166; 
wire N167; 
wire N168; 
wire N169; 
wire N170; 
wire N171; 
wire N172; 
wire N173; 
wire N174; 
wire N175; 
wire N176; 
wire N177; 
wire N178; 
wire N179; 
wire N180; 
wire N181; 
wire N182; 
wire N183; 
wire N184; 
wire N185; 
wire N186; 
wire N187; 
wire N188; 
wire N189; 
wire N190; 
wire N191; 
wire N192; 
wire N193; 
wire N194; 
wire N195; 
wire N196; 
wire N197; 
wire N198; 
wire N199; 
wire N200; 
wire N201; 
wire N202; 
wire N203; 
wire N204; 
wire N205; 
wire N206; 
wire N207; 
wire N208; 
wire N209; 
wire N210; 
wire N211; 
wire N212; 
wire N213; 
wire N214; 
wire N215; 
wire N216; 
wire N217; 
wire N218; 
wire N219; 
wire N220; 
wire N221; 
wire N222; 
wire N223; 
wire N224; 
wire N225; 
wire N226; 
wire N227; 
wire N228; 
wire N229; 
wire N230; 
wire N231; 
wire N232; 
wire N233; 
wire N234; 
wire N235; 
wire N236; 
wire N237; 
wire N238; 
wire N239; 
wire N240; 
wire N241; 
wire N242; 
wire N243; 
wire N244; 
wire N245; 
wire N246; 
wire N247; 
wire N248; 
wire N249; 
wire N250; 
wire N251; 
wire N252; 
wire N253; 
wire N254; 
wire N255; 
wire N256; 
wire N257; 
wire N258; 
wire N259; 
wire N260; 
wire N261; 
wire N262; 
wire N263; 
wire N264; 
wire N265; 
wire N266; 
wire N267; 
wire N268; 
wire N269; 
wire N270; 
wire N271; 
wire N272; 
wire N273; 
wire N274; 
wire N275; 
wire N276; 
wire N277; 
wire N278; 
wire N279; 
wire N280; 
wire N281; 
wire N282; 
wire N283; 
wire N284; 
wire N285; 
wire N286; 
wire N287; 
wire N288; 
wire N289; 
wire N290; 
wire N291; 
wire N292; 
wire N293; 
wire N294; 
wire N295; 
wire N296; 
wire N297; 
wire N298; 
wire N299; 
wire N300; 
wire N301; 
wire N302; 
wire N303; 
wire N304; 
wire N305; 
wire N306; 
wire N307; 
wire N308; 
wire N309; 
wire N310; 
wire N311; 
wire N312; 
wire N313; 
wire N314; 
wire N315; 
wire N316; 
wire N317; 
wire N318; 
wire N319; 
wire N320; 
wire N321; 
wire N322; 
wire N323; 
wire N324; 
wire N325; 
wire N326; 
wire N327; 
wire N328; 
wire N329; 
wire N330; 
wire N331; 
wire N332; 
wire N333; 
wire N334; 
wire N335; 
wire N336; 
wire N337; 
wire N338; 
wire N339; 
wire N340; 
wire N341; 
wire N342; 
wire N343; 
wire N344; 
wire N345; 
wire N346; 
wire N347; 
wire N348; 
wire N349; 
wire N350; 
wire N351; 
wire N352; 
wire N353; 
wire N354; 
wire N355; 
wire N356; 
wire N357; 
wire N358; 
wire N359; 
wire N360; 
wire N361; 
wire N362; 
wire N363; 
wire N364; 
wire N365; 
wire N366; 
wire N367; 
wire N368; 
wire N369; 
wire N370; 
wire N371; 
wire N372; 
wire N373; 
wire N374; 
wire N375; 
wire N376; 
wire N377; 
wire N378; 
wire N379; 
wire N380; 
wire N381; 
wire N382; 
wire N383; 
wire N384; 
wire N385; 
wire N386; 
wire N387; 
wire N388; 
wire N389; 
wire N390; 
wire N391; 
wire N392; 
wire N393; 
wire N394; 
wire N395; 
wire N396; 
wire N397; 
wire N398; 
wire N399; 
wire N400; 
wire N401; 
wire N402; 
wire N403; 
wire N404; 
wire N405; 
wire N406; 
wire N407; 
wire N408; 
wire N409; 
wire N410; 
wire N411; 
wire N412; 
wire N413; 
wire N414; 
wire N415; 
wire N416; 
wire N417; 
wire N418; 
wire N419; 
wire N420; 
wire N421; 
wire N422; 
wire N423; 
wire N424; 
wire N425; 
wire N426; 
wire N427; 
wire N428; 
wire N429; 
wire N430; 
wire N431; 
wire N432; 
wire N433; 
wire N434; 
wire N435; 
wire N436; 
wire N437; 
wire N438; 
wire N439; 
wire N440; 
wire N441; 
wire N442; 
wire N443; 
wire N444; 

assign N14 = ~(N7); 
assign N15 = ~(N3); 
assign N16 = N8 & N2; 
assign N17 = ~(N1); 
assign N18 = ~(N7); 
assign N19 = ~(N11); 
assign N20 = ~(N5); 
assign N21 = ~(N4); 
assign N22 = ~(N1); 
assign N23 = ~(N4); 
assign N24 = ~(N10); 
assign N25 = ~(N8); 
assign N26 = ~(N6); 
assign N27 = ~(N2); 
assign N28 = ~(N7); 
assign N29 = ~(N3); 
assign N30 = ~(N6); 
assign N31 = ~(N30); 
assign N32 = ~(N13); 
assign N33 = ~(N14); 
assign N34 = ~(N1); 
assign N35 = ~(N21); 
assign N36 = N26 & N4; 
assign N37 = ~(N6); 
assign N38 = ~(N7); 
assign N39 = ~(N21); 
assign N40 = ~(N1); 
assign N41 = ~(N26); 
assign N42 = ~(N3); 
assign N43 = ~(N24); 
assign N44 = ~(N11); 
assign N45 = ~(N21); 
assign N46 = ~(N9); 
assign N47 = ~(N26); 
assign N48 = N13 & N22 & N15; 
assign N49 = ~(N12); 
assign N50 = ~(N15); 
assign N51 = ~(N14); 
assign N52 = ~(N23); 
assign N53 = ~(N2); 
assign N54 = N6 | N3; 
assign N55 = ~(N18); 
assign N56 = ~(N24); 
assign N57 = ~(N9); 
assign N58 = ~(N21); 
assign N59 = N27 & N28 & N20; 
assign N60 = N20 | N22; 
assign N61 = ~(N22); 
assign N62 = ~(N48); 
assign N63 = N25 & N49; 
assign N64 = ~(N6); 
assign N65 = N17 & N32; 
assign N66 = ~(N5); 
assign N67 = ~(N5); 
assign N68 = ~(N2); 
assign N69 = ~(N24); 
assign N70 = N48 & N60; 
assign N71 = N24 | N57 | N59; 
assign N72 = N63 | N46; 
assign N73 = N30 & N61; 
assign N74 = N52 | N63; 
assign N75 = N51 | N23; 
assign N76 = ~(N16); 
assign N77 = ~(N73); 
assign N78 = ~(N69); 
assign N79 = ~(N57); 
assign N80 = ~(N58); 
assign N81 = ~(N53); 
assign N82 = ~(N20); 
assign N83 = ~(N68); 
assign N84 = ~(N19); 
assign N85 = ~(N56); 
assign N86 = ~(N54); 
assign N87 = ~(N66); 
assign N88 = ~(N11); 
assign N89 = ~(N75); 
assign N90 = ~(N25); 
assign N91 = ~(N51); 
assign N92 = ~(N5); 
assign N93 = ~(N71); 
assign N94 = ~(N18); 
assign N95 = ~(N54); 
assign N96 = ~(N25); 
assign N97 = ~(N11); 
assign N98 = ~(N41); 
assign N99 = N49 | N70; 
assign N100 = ~(N3); 
assign N101 = N71 | N69; 
assign N102 = ~(N70); 
assign N103 = ~(N74); 
assign N104 = N14 | N15; 
assign N105 = ~(N45); 
assign N106 = ~(N75); 
assign N107 = ~(N54); 
assign N108 = ~(N59); 
assign N109 = ~(N72); 
assign N110 = ~(N25); 
assign N111 = ~(N70); 
assign N112 = ~(N11); 
assign N113 = ~(N25); 
assign N114 = ~(N36); 
assign N115 = ~(N50); 
assign N116 = ~(N56); 
assign N117 = ~(N75); 
assign N118 = ~(N75); 
assign N119 = ~(N53); 
assign N120 = ~(N70); 
assign N121 = ~(N41); 
assign N122 = ~(N36); 
assign N123 = ~(N60); 
assign N124 = N33 & N52; 
assign N125 = ~(N19); 
assign N126 = ~(N66); 
assign N127 = ~(N58); 
assign N128 = ~(N35); 
assign N129 = ~(N4); 
assign N130 = ~(N124); 
assign N131 = ~(N73); 
assign N132 = ~(N30); 
assign N133 = ~(N29); 
assign N134 = ~(N36); 
assign N135 = ~(N97); 
assign N136 = ~(N50); 
assign N137 = ~(N61); 
assign N138 = ~(N57); 
assign N139 = ~(N41); 
assign N140 = ~(N12); 
assign N141 = ~(N10); 
assign N142 = ~(N105); 
assign N143 = ~(N39); 
assign N144 = ~(N16); 
assign N145 = ~(N57); 
assign N146 = ~(N39); 
assign N147 = ~(N56); 
assign N148 = ~(N70); 
assign N149 = N19 & N75; 
assign N150 = ~(N72); 
assign N151 = ~(N43); 
assign N152 = ~(N23); 
assign N153 = ~(N73); 
assign N154 = ~(N72); 
assign N155 = N73 & N60; 
assign N156 = ~(N59); 
assign N157 = ~(N60); 
assign N158 = N78 & N65; 
assign N159 = ~(N96); 
assign N160 = ~(N73); 
assign N161 = ~(N50); 
assign N162 = N106 & N74; 
assign N163 = ~(N116); 
assign N164 = ~(N29); 
assign N165 = N114 | N73; 
assign N166 = ~(N109); 
assign N167 = ~(N65); 
assign N168 = ~(N48); 
assign N169 = N95 & N12; 
assign N170 = ~(N41); 
assign N171 = N121 & N92; 
assign N172 = N119 | N22; 
assign N173 = ~(N24); 
assign N174 = ~(N10); 
assign N175 = ~(N112); 
assign N176 = ~(N71); 
assign N177 = ~(N12); 
assign N178 = ~(N63); 
assign N179 = ~(N42); 
assign N180 = ~(N50); 
assign N181 = N62 & N61; 
assign N182 = ~(N37); 
assign N183 = ~(N150); 
assign N184 = ~(N71); 
assign N185 = ~(N14); 
assign N186 = ~(N74); 
assign N187 = N108 | N43; 
assign N188 = ~(N57); 
assign N189 = ~(N17); 
assign N190 = ~(N26); 
assign N191 = ~(N46); 
assign N192 = N23 & N9; 
assign N193 = ~(N107); 
assign N194 = ~(N174); 
assign N195 = ~(N65); 
assign N196 = ~(N140); 
assign N197 = ~(N82); 
assign N198 = ~(N37); 
assign N199 = N118 & N54; 
assign N200 = ~(N53); 
assign N201 = ~(N112); 
assign N202 = N12 | N71; 
assign N203 = N169 & N168; 
assign N204 = ~(N112); 
assign N205 = N43 & N141; 
assign N206 = ~(N58); 
assign N207 = ~(N156); 
assign N208 = N46 & N61 & N94; 
assign N209 = ~(N120); 
assign N210 = ~(N151); 
assign N211 = ~(N150); 
assign N212 = ~(N162); 
assign N213 = ~(N55); 
assign N214 = ~(N96); 
assign N215 = ~(N9); 
assign N216 = ~(N15); 
assign N217 = ~(N47); 
assign N218 = N4 & N167 & N65; 
assign N219 = N133 & N172; 
assign N220 = ~(N102); 
assign N221 = ~(N93); 
assign N222 = N120 & N118; 
assign N223 = N102 & N74; 
assign N224 = ~(N217); 
assign N225 = ~(N154); 
assign N226 = N1 | N141; 
assign N227 = ~(N145); 
assign N228 = N81 | N44; 
assign N229 = N147 | N16; 
assign N230 = N122 | N68; 
assign N231 = N82 & N118; 
assign N232 = ~(N183); 
assign N233 = N192 & N101; 
assign N234 = ~(N177); 
assign N235 = ~(N87); 
assign N236 = ~(N17); 
assign N237 = ~(N58); 
assign N238 = N70 | N143; 
assign N239 = ~(N44); 
assign N240 = ~(N151); 
assign N241 = N162 & N182; 
assign N242 = ~(N155); 
assign N243 = ~(N74); 
assign N244 = N180 & N196 & N211 & N66; 
assign N245 = ~(N165); 
assign N246 = ~(N175); 
assign N247 = N148 & N134; 
assign N248 = ~(N181); 
assign N249 = N123 | N152; 
assign N250 = ~(N68); 
assign N251 = ~(N39); 
assign N252 = N38 | N63; 
assign N253 = N16 & N213; 
assign N254 = ~(N184); 
assign N255 = ~(N85); 
assign N256 = ~(N195); 
assign N257 = ~(N214); 
assign N258 = ~(N16); 
assign N259 = N190 & N55; 
assign N260 = ~(N23); 
assign N261 = ~(N118); 
assign N262 = ~(N39); 
assign N263 = ~(N67); 
assign N264 = ~(N26); 
assign N265 = ~(N20); 
assign N266 = N250 & N195; 
assign N267 = N64 | N80; 
assign N268 = ~(N129); 
assign N269 = ~(N145); 
assign N270 = ~(N103); 
assign N271 = ~(N102); 
assign N272 = N157 | N196; 
assign N273 = ~(N8); 
assign N274 = N2 & N101; 
assign N275 = ~(N82); 
assign N276 = ~(N182); 
assign N277 = N185 | N224; 
assign N278 = ~(N190); 
assign N279 = N237 & N44; 
assign N280 = ~(N108); 
assign N281 = ~(N69); 
assign N282 = N131 & N28; 
assign N283 = ~(N193); 
assign N284 = ~(N172); 
assign N285 = N29 & N188; 
assign N286 = ~(N63); 
assign N287 = ~(N81); 
assign N288 = N67 & N180; 
assign N289 = ~(N196); 
assign N290 = ~(N14); 
assign N291 = N11 & N26; 
assign N292 = ~(N248); 
assign N293 = ~(N43); 
assign N294 = ~(N196); 
assign N295 = ~(N221); 
assign N296 = ~(N156); 
assign N297 = ~(N119); 
assign N298 = N79 & N66; 
assign N299 = ~(N96); 
assign N300 = ~(N66); 
assign N301 = ~(N134); 
assign N302 = ~(N5); 
assign N303 = N239 & N148; 
assign N304 = ~(N202); 
assign N305 = ~(N171); 
assign N306 = N168 | N213 | N247; 
assign N307 = N205 & N220 & N87; 
assign N308 = ~(N197); 
assign N309 = N142 & N195; 
assign N310 = N155 & N240; 
assign N311 = ~(N63); 
assign N312 = ~(N100); 
assign N313 = ~(N52); 
assign N314 = ~(N55); 
assign N315 = N174 | N129; 
assign N316 = ~(N8); 
assign N317 = N56 & N8; 
assign N318 = N187 & N216 & N92; 
assign N319 = ~(N19); 
assign N320 = N21 & N60 & N202 & N22; 
assign N321 = N197 & N304 & N61; 
assign N322 = N50 | N207; 
assign N323 = N41 & N288; 
assign N324 = N77 | N103 | N236 | N124; 
assign N325 = N231 & N13; 
assign N326 = N10 & N243 & N263 & N72; 
assign N327 = ~(N159); 
assign N328 = N40 & N153 & N213; 
assign N329 = N271 | N145; 
assign N330 = ~(N229); 
assign N331 = ~(N249); 
assign N332 = N107 & N194; 
assign N333 = N92 | N176 | N245 | N260 | N296 | N178; 
assign N334 = N138 | N229 | N308; 
assign N335 = N132 | N312 | N209; 
assign N336 = N127 & N284 & N288; 
assign N337 = N7 | N34 | N55 | N223 | N238 | N242 | N256 | N186; 
assign N338 = N143 & N179 & N254 & N272 & N282; 
assign N339 = N99 & N183 & N189 & N323 & N152; 
assign N340 = N164 | N170 | N314 | N318; 
assign N341 = N156 | N104; 
assign N342 = N9 & N109 & N218 & N16; 
assign N343 = N232 | N326 | N283 | N275; 
assign N344 = N15 & N306; 
assign N345 = N85 | N96 | N68; 
assign N346 = N199 | N251 | N280 | N179; 
assign N347 = N47 | N86 | N129 | N209 | N226 | N123; 
assign N348 = N45 & N91 & N191 & N266 & N329; 
assign N349 = ~(N121); 
assign N350 = N39 | N234 | N253 | N277 | N283 | N287 | N298 | N310; 
assign N351 = N32 | N100 | N336 | N337; 
assign N352 = N35 & N36 & N44 & N65 & N68 & N140 & N188 & N235; 
assign N353 = N88 & N116 & N204 & N315 & N340 & N346 & N135; 
assign N354 = N18 & N37 & N54 & N177 & N208 & N210 & N259 & N297; 
assign N355 = N125 | N326; 
assign N356 = N160 | N181 | N247; 
assign N357 = N75 & N137 & N317 & N351 & N254; 
assign N358 = ~(N61); 
assign N359 = N31 | N227 | N255 | N343 | N234; 
assign N360 = N130 & N233 & N59; 
assign N361 = ~(N319); 
assign N362 = ~(N244); 
assign N363 = ~(N315); 
assign N364 = ~(N233); 
assign N365 = N83 | N184 | N273 | N305; 
assign N366 = N139 & N206 & N228 & N258 & N290; 
assign N367 = N90 & N135 & N172 & N269 & N281; 
assign N368 = N215 | N219 | N345 | N163; 
assign N369 = N84 & N248; 
assign N370 = N173 & N198; 
assign N371 = N311 | N17; 
assign N372 = N98 | N333 | N207; 
assign N373 = N105 | N146 | N35; 
assign N374 = ~(N283); 
assign N375 = N69 | N188; 
assign N376 = ~(N178); 
assign N377 = N203 | N262 | N356 | N230; 
assign N378 = N330 | N234; 
assign N379 = N257 | N289 | N348 | N313; 
assign N380 = ~(N13); 
assign N381 = ~(N58); 
assign N382 = N294 | N119; 
assign N383 = N358 | N224; 
assign N384 = ~(N68); 
assign N385 = ~(N241); 
assign N386 = N113 | N217 | N352 | N112; 
assign N387 = ~(N13); 
assign N388 = N165 | N316 | N256; 
assign N389 = ~(N250); 
assign N390 = N93 | N121; 
assign N391 = ~(N43); 
assign N392 = N126 | N254; 
assign N393 = ~(N318); 
assign N394 = N128 | N246 | N335 | N338 | N62; 
assign N395 = N72 | N117 | N225; 
assign N396 = ~(N126); 
assign N397 = N362 | N19 | N292; 
assign N398 = N193 & N249 & N303 & N328; 
assign N399 = N279 & N359 & N235; 
assign N400 = N186 | N108; 
assign N401 = ~(N296); 
assign N402 = N136 & N175 & N285 & N145; 
assign N403 = ~(N249); 
assign N404 = ~(N347); 
assign N405 = ~(N350); 
assign N406 = N274 | N309 | N318 | N344 | N365 | N321; 
assign N407 = N295 & N369 & N375 & N259; 
assign N408 = N178 & N382; 
assign N409 = N149 & N163; 
assign N410 = ~(N59); 
assign N411 = ~(N62); 
assign N412 = N319 & N250; 
assign N413 = N322 & N389; 
assign N414 = ~(N256); 
assign N415 = ~(N103); 
assign N416 = N201 | N252 | N391 | N175; 
assign N417 = ~(N403); 
assign N418 = N307 & N320 & N355 & N363 & N76; 
assign N419 = N258 & N394; 
assign N420 = N261 & N327 & N373 & N388 & N123; 
assign N421 = N110 | N160; 
assign N422 = N377 & N78 & N347; 
assign N423 = N276 & N368 & N319; 
assign N424 = N396 | N62; 
assign N425 = N145 & N197; 
assign N426 = N291 | N386 | N148; 
assign N427 = N384 & N402; 
assign N428 = N154 | N171 | N122; 
assign N429 = N144 | N158 | N264 | N69; 
assign N430 = N395 & N155; 
assign N431 = ~(N215); 
assign N432 = N286 | N379 | N306; 
assign N433 = N161 | N300 | N147; 
assign N434 = ~(N231); 
assign N435 = N282 & N361 & N178; 
assign N436 = N399 & N195; 
assign N437 = N331 & N154; 
assign N438 = N378 | N139; 
assign N439 = ~(N333); 
assign N440 = ~(N180); 
assign N441 = ~(N278); 
assign N442 = ~(N195); 
assign N443 = N383 & N387 & N121; 
assign N444 = N404 & N218; 
assign N445 = N166 | N354 | N429 | N440; 
assign N446 = ~(N360); 
assign N447 = N299 & N357 & N364 & N408 & N426 & N434; 
assign N448 = N265 | N270 | N353 | N418; 
assign N449 = N400 | N406 | N435; 
assign N450 = N76 | N302 | N405; 
assign N451 = N367 | N370 | N393; 
assign N452 = ~(N145); 
assign N453 = N332 | N409 | N420 | N421 | N425; 
assign N454 = N417 | N442 | N444; 
assign N455 = N313 | N392 | N407 | N415 | N424; 
assign N456 = N115 & N247; 
assign N457 = N224 | N374 | N433; 
assign N458 = N124 & N230 & N293 & N381 & N413 & N414 & N416 & N427; 
assign N459 = N101 & N366 & N385; 
assign N460 = N268 & N390 & N428; 
assign N461 = N111 | N221 | N401 | N422 | N430 | N441; 
assign N462 = ~(N200); 
assign N463 = N324 & N341 & N431 & N437; 
assign N464 = N152 & N212 & N301 & N397 & N436; 
assign N465 = N207 & N398 & N432; 
assign N466 = N89 | N410; 
assign N467 = N339 | N376 | N411; 
assign N468 = ~(N371); 
assign N469 = N104 & N267 & N372 & N380; 
assign N470 = N225 & N325 & N412 & N419 & N423 & N439 & N342 & N443; 
assign N471 = N222 & N334 & N349 & N438; 
endmodule
