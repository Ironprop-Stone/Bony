module Depth_10_20_Nodes_200_400_S004 (N1, N2, N3, N4, N5, N318, N319, N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330, N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341, N342);

input N1; 
input N2; 
input N3; 
input N4; 
input N5; 

output N318; 
output N319; 
output N320; 
output N321; 
output N322; 
output N323; 
output N324; 
output N325; 
output N326; 
output N327; 
output N328; 
output N329; 
output N330; 
output N331; 
output N332; 
output N333; 
output N334; 
output N335; 
output N336; 
output N337; 
output N338; 
output N339; 
output N340; 
output N341; 
output N342; 

wire N6; 
wire N7; 
wire N8; 
wire N9; 
wire N10; 
wire N11; 
wire N12; 
wire N13; 
wire N14; 
wire N15; 
wire N16; 
wire N17; 
wire N18; 
wire N19; 
wire N20; 
wire N21; 
wire N22; 
wire N23; 
wire N24; 
wire N25; 
wire N26; 
wire N27; 
wire N28; 
wire N29; 
wire N30; 
wire N31; 
wire N32; 
wire N33; 
wire N34; 
wire N35; 
wire N36; 
wire N37; 
wire N38; 
wire N39; 
wire N40; 
wire N41; 
wire N42; 
wire N43; 
wire N44; 
wire N45; 
wire N46; 
wire N47; 
wire N48; 
wire N49; 
wire N50; 
wire N51; 
wire N52; 
wire N53; 
wire N54; 
wire N55; 
wire N56; 
wire N57; 
wire N58; 
wire N59; 
wire N60; 
wire N61; 
wire N62; 
wire N63; 
wire N64; 
wire N65; 
wire N66; 
wire N67; 
wire N68; 
wire N69; 
wire N70; 
wire N71; 
wire N72; 
wire N73; 
wire N74; 
wire N75; 
wire N76; 
wire N77; 
wire N78; 
wire N79; 
wire N80; 
wire N81; 
wire N82; 
wire N83; 
wire N84; 
wire N85; 
wire N86; 
wire N87; 
wire N88; 
wire N89; 
wire N90; 
wire N91; 
wire N92; 
wire N93; 
wire N94; 
wire N95; 
wire N96; 
wire N97; 
wire N98; 
wire N99; 
wire N100; 
wire N101; 
wire N102; 
wire N103; 
wire N104; 
wire N105; 
wire N106; 
wire N107; 
wire N108; 
wire N109; 
wire N110; 
wire N111; 
wire N112; 
wire N113; 
wire N114; 
wire N115; 
wire N116; 
wire N117; 
wire N118; 
wire N119; 
wire N120; 
wire N121; 
wire N122; 
wire N123; 
wire N124; 
wire N125; 
wire N126; 
wire N127; 
wire N128; 
wire N129; 
wire N130; 
wire N131; 
wire N132; 
wire N133; 
wire N134; 
wire N135; 
wire N136; 
wire N137; 
wire N138; 
wire N139; 
wire N140; 
wire N141; 
wire N142; 
wire N143; 
wire N144; 
wire N145; 
wire N146; 
wire N147; 
wire N148; 
wire N149; 
wire N150; 
wire N151; 
wire N152; 
wire N153; 
wire N154; 
wire N155; 
wire N156; 
wire N157; 
wire N158; 
wire N159; 
wire N160; 
wire N161; 
wire N162; 
wire N163; 
wire N164; 
wire N165; 
wire N166; 
wire N167; 
wire N168; 
wire N169; 
wire N170; 
wire N171; 
wire N172; 
wire N173; 
wire N174; 
wire N175; 
wire N176; 
wire N177; 
wire N178; 
wire N179; 
wire N180; 
wire N181; 
wire N182; 
wire N183; 
wire N184; 
wire N185; 
wire N186; 
wire N187; 
wire N188; 
wire N189; 
wire N190; 
wire N191; 
wire N192; 
wire N193; 
wire N194; 
wire N195; 
wire N196; 
wire N197; 
wire N198; 
wire N199; 
wire N200; 
wire N201; 
wire N202; 
wire N203; 
wire N204; 
wire N205; 
wire N206; 
wire N207; 
wire N208; 
wire N209; 
wire N210; 
wire N211; 
wire N212; 
wire N213; 
wire N214; 
wire N215; 
wire N216; 
wire N217; 
wire N218; 
wire N219; 
wire N220; 
wire N221; 
wire N222; 
wire N223; 
wire N224; 
wire N225; 
wire N226; 
wire N227; 
wire N228; 
wire N229; 
wire N230; 
wire N231; 
wire N232; 
wire N233; 
wire N234; 
wire N235; 
wire N236; 
wire N237; 
wire N238; 
wire N239; 
wire N240; 
wire N241; 
wire N242; 
wire N243; 
wire N244; 
wire N245; 
wire N246; 
wire N247; 
wire N248; 
wire N249; 
wire N250; 
wire N251; 
wire N252; 
wire N253; 
wire N254; 
wire N255; 
wire N256; 
wire N257; 
wire N258; 
wire N259; 
wire N260; 
wire N261; 
wire N262; 
wire N263; 
wire N264; 
wire N265; 
wire N266; 
wire N267; 
wire N268; 
wire N269; 
wire N270; 
wire N271; 
wire N272; 
wire N273; 
wire N274; 
wire N275; 
wire N276; 
wire N277; 
wire N278; 
wire N279; 
wire N280; 
wire N281; 
wire N282; 
wire N283; 
wire N284; 
wire N285; 
wire N286; 
wire N287; 
wire N288; 
wire N289; 
wire N290; 
wire N291; 
wire N292; 
wire N293; 
wire N294; 
wire N295; 
wire N296; 
wire N297; 
wire N298; 
wire N299; 
wire N300; 
wire N301; 
wire N302; 
wire N303; 
wire N304; 
wire N305; 
wire N306; 
wire N307; 
wire N308; 
wire N309; 
wire N310; 
wire N311; 
wire N312; 
wire N313; 
wire N314; 
wire N315; 
wire N316; 
wire N317; 

assign N6 = ~(N5); 
assign N7 = N5 & N1; 
assign N8 = ~(N1); 
assign N9 = ~(N2); 
assign N10 = ~(N5); 
assign N11 = ~(N3); 
assign N12 = ~(N1); 
assign N13 = ~(N2); 
assign N14 = ~(N2); 
assign N15 = ~(N1); 
assign N16 = ~(N5); 
assign N17 = ~(N5); 
assign N18 = ~(N12); 
assign N19 = ~(N1); 
assign N20 = ~(N3); 
assign N21 = ~(N10); 
assign N22 = ~(N10); 
assign N23 = ~(N4); 
assign N24 = ~(N11); 
assign N25 = N8 & N11; 
assign N26 = ~(N2); 
assign N27 = N6 & N15; 
assign N28 = ~(N9); 
assign N29 = ~(N16); 
assign N30 = ~(N10); 
assign N31 = ~(N17); 
assign N32 = ~(N9); 
assign N33 = ~(N4); 
assign N34 = ~(N3); 
assign N35 = ~(N4); 
assign N36 = ~(N11); 
assign N37 = ~(N6); 
assign N38 = ~(N10); 
assign N39 = ~(N7); 
assign N40 = ~(N11); 
assign N41 = ~(N16); 
assign N42 = ~(N14); 
assign N43 = ~(N6); 
assign N44 = ~(N16); 
assign N45 = ~(N11); 
assign N46 = ~(N7); 
assign N47 = ~(N16); 
assign N48 = ~(N8); 
assign N49 = ~(N17); 
assign N50 = ~(N15); 
assign N51 = ~(N4); 
assign N52 = ~(N15); 
assign N53 = ~(N4); 
assign N54 = ~(N14); 
assign N55 = ~(N17); 
assign N56 = ~(N2); 
assign N57 = ~(N7); 
assign N58 = ~(N5); 
assign N59 = ~(N8); 
assign N60 = ~(N17); 
assign N61 = ~(N12); 
assign N62 = ~(N56); 
assign N63 = ~(N44); 
assign N64 = N29 & N14; 
assign N65 = N21 & N8; 
assign N66 = ~(N41); 
assign N67 = ~(N20); 
assign N68 = ~(N27); 
assign N69 = ~(N3); 
assign N70 = ~(N7); 
assign N71 = ~(N41); 
assign N72 = ~(N17); 
assign N73 = ~(N15); 
assign N74 = ~(N21); 
assign N75 = ~(N10); 
assign N76 = ~(N47); 
assign N77 = N53 | N56 | N27; 
assign N78 = N58 & N26; 
assign N79 = ~(N53); 
assign N80 = ~(N38); 
assign N81 = ~(N13); 
assign N82 = ~(N15); 
assign N83 = ~(N51); 
assign N84 = ~(N53); 
assign N85 = ~(N29); 
assign N86 = N38 | N16; 
assign N87 = N49 | N36; 
assign N88 = ~(N15); 
assign N89 = N16 & N12; 
assign N90 = ~(N31); 
assign N91 = ~(N35); 
assign N92 = N37 & N9; 
assign N93 = ~(N29); 
assign N94 = ~(N38); 
assign N95 = N48 & N12; 
assign N96 = ~(N9); 
assign N97 = ~(N40); 
assign N98 = ~(N3); 
assign N99 = ~(N56); 
assign N100 = N3 | N27; 
assign N101 = ~(N98); 
assign N102 = ~(N62); 
assign N103 = N97 | N55; 
assign N104 = N71 & N25; 
assign N105 = ~(N87); 
assign N106 = N92 | N39; 
assign N107 = ~(N55); 
assign N108 = ~(N39); 
assign N109 = N77 | N22; 
assign N110 = ~(N76); 
assign N111 = ~(N65); 
assign N112 = N52 & N79 & N62; 
assign N113 = ~(N44); 
assign N114 = ~(N8); 
assign N115 = ~(N25); 
assign N116 = N42 & N68; 
assign N117 = N17 & N47; 
assign N118 = ~(N29); 
assign N119 = ~(N66); 
assign N120 = N68 | N9; 
assign N121 = ~(N14); 
assign N122 = ~(N62); 
assign N123 = ~(N20); 
assign N124 = ~(N99); 
assign N125 = N72 | N55; 
assign N126 = ~(N86); 
assign N127 = ~(N99); 
assign N128 = ~(N88); 
assign N129 = ~(N44); 
assign N130 = ~(N26); 
assign N131 = N40 | N70; 
assign N132 = ~(N50); 
assign N133 = ~(N61); 
assign N134 = N73 | N76; 
assign N135 = ~(N129); 
assign N136 = ~(N107); 
assign N137 = ~(N92); 
assign N138 = ~(N108); 
assign N139 = ~(N112); 
assign N140 = N13 & N106; 
assign N141 = N86 | N67; 
assign N142 = ~(N76); 
assign N143 = N100 | N79; 
assign N144 = N2 | N121 | N142; 
assign N145 = ~(N84); 
assign N146 = ~(N108); 
assign N147 = ~(N84); 
assign N148 = N103 & N82; 
assign N149 = ~(N79); 
assign N150 = ~(N8); 
assign N151 = ~(N6); 
assign N152 = ~(N65); 
assign N153 = ~(N20); 
assign N154 = ~(N97); 
assign N155 = ~(N78); 
assign N156 = ~(N128); 
assign N157 = N132 & N143; 
assign N158 = ~(N30); 
assign N159 = ~(N26); 
assign N160 = N118 & N71; 
assign N161 = ~(N143); 
assign N162 = ~(N13); 
assign N163 = ~(N107); 
assign N164 = ~(N13); 
assign N165 = ~(N83); 
assign N166 = ~(N22); 
assign N167 = ~(N34); 
assign N168 = ~(N117); 
assign N169 = N119 & N109; 
assign N170 = ~(N106); 
assign N171 = ~(N6); 
assign N172 = ~(N112); 
assign N173 = N66 | N71; 
assign N174 = ~(N23); 
assign N175 = ~(N92); 
assign N176 = ~(N90); 
assign N177 = ~(N47); 
assign N178 = ~(N133); 
assign N179 = ~(N81); 
assign N180 = ~(N63); 
assign N181 = ~(N107); 
assign N182 = ~(N141); 
assign N183 = ~(N69); 
assign N184 = ~(N81); 
assign N185 = ~(N36); 
assign N186 = ~(N73); 
assign N187 = ~(N12); 
assign N188 = ~(N68); 
assign N189 = ~(N87); 
assign N190 = ~(N107); 
assign N191 = ~(N34); 
assign N192 = ~(N25); 
assign N193 = ~(N36); 
assign N194 = ~(N73); 
assign N195 = N23 & N82 & N112; 
assign N196 = ~(N140); 
assign N197 = ~(N122); 
assign N198 = N101 & N126; 
assign N199 = ~(N89); 
assign N200 = ~(N32); 
assign N201 = ~(N129); 
assign N202 = ~(N120); 
assign N203 = ~(N143); 
assign N204 = N1 & N52; 
assign N205 = ~(N36); 
assign N206 = ~(N63); 
assign N207 = ~(N27); 
assign N208 = ~(N94); 
assign N209 = N115 & N90; 
assign N210 = ~(N38); 
assign N211 = ~(N134); 
assign N212 = N25 | N98; 
assign N213 = ~(N46); 
assign N214 = ~(N108); 
assign N215 = N30 | N124; 
assign N216 = N12 & N34; 
assign N217 = ~(N129); 
assign N218 = ~(N122); 
assign N219 = ~(N98); 
assign N220 = ~(N142); 
assign N221 = N11 & N40; 
assign N222 = ~(N13); 
assign N223 = ~(N23); 
assign N224 = ~(N107); 
assign N225 = ~(N125); 
assign N226 = ~(N109); 
assign N227 = ~(N132); 
assign N228 = ~(N69); 
assign N229 = ~(N41); 
assign N230 = ~(N85); 
assign N231 = ~(N138); 
assign N232 = ~(N131); 
assign N233 = ~(N33); 
assign N234 = ~(N120); 
assign N235 = ~(N89); 
assign N236 = ~(N137); 
assign N237 = ~(N18); 
assign N238 = N80 | N128 | N168 | N204 | N25; 
assign N239 = ~(N112); 
assign N240 = ~(N46); 
assign N241 = ~(N129); 
assign N242 = ~(N124); 
assign N243 = ~(N158); 
assign N244 = ~(N230); 
assign N245 = ~(N106); 
assign N246 = ~(N120); 
assign N247 = ~(N115); 
assign N248 = N4 & N93 & N33; 
assign N249 = ~(N131); 
assign N250 = N55 & N231; 
assign N251 = ~(N162); 
assign N252 = ~(N222); 
assign N253 = ~(N129); 
assign N254 = N45 & N234 & N135; 
assign N255 = ~(N231); 
assign N256 = ~(N198); 
assign N257 = ~(N178); 
assign N258 = N159 | N211 | N235; 
assign N259 = N193 & N14; 
assign N260 = ~(N190); 
assign N261 = ~(N40); 
assign N262 = N18 | N139; 
assign N263 = ~(N74); 
assign N264 = ~(N40); 
assign N265 = N176 | N220 | N138; 
assign N266 = N135 & N197 & N233; 
assign N267 = N61 | N136; 
assign N268 = ~(N214); 
assign N269 = ~(N34); 
assign N270 = ~(N92); 
assign N271 = ~(N107); 
assign N272 = ~(N110); 
assign N273 = N96 | N130; 
assign N274 = ~(N133); 
assign N275 = ~(N206); 
assign N276 = ~(N138); 
assign N277 = ~(N138); 
assign N278 = ~(N132); 
assign N279 = ~(N47); 
assign N280 = N156 | N39; 
assign N281 = ~(N137); 
assign N282 = ~(N146); 
assign N283 = N41 & N111 & N143; 
assign N284 = N46 | N140; 
assign N285 = N198 | N202 | N113; 
assign N286 = N84 | N194 | N133; 
assign N287 = ~(N224); 
assign N288 = N109 & N158; 
assign N289 = N218 & N132; 
assign N290 = ~(N215); 
assign N291 = N14 | N210 | N68; 
assign N292 = N91 | N178; 
assign N293 = ~(N131); 
assign N294 = ~(N201); 
assign N295 = N19 & N31 & N114 & N153 & N186 & N232 & N40; 
assign N296 = N57 & N78 & N127 & N196 & N252 & N283; 
assign N297 = N141 | N157 | N224 | N292 | N282; 
assign N298 = N81 | N136 | N212 | N142 | N291; 
assign N299 = N122 & N130 & N167 & N200 & N221 & N270 & N281 & N121; 
assign N300 = N10 & N146 & N177 & N205 & N229 & N256 & N271 & N273; 
assign N301 = N182 | N233 | N244 | N277 | N255; 
assign N302 = N28 & N187 & N226 & N242 & N55; 
assign N303 = N32 | N85 | N192 | N138; 
assign N304 = N216 | N217 | N219 | N92; 
assign N305 = N54 & N69 & N74 & N140 & N171 & N209 & N245 & N261; 
assign N306 = N44 & N102 & N113 & N123 & N124 & N145 & N165 & N222; 
assign N307 = N161 & N175 & N183 & N185; 
assign N308 = N27 | N138 | N163 | N188 | N180; 
assign N309 = N120 | N228; 
assign N310 = N36 | N75 | N87 | N131 | N133 | N259 | N280 | N300; 
assign N311 = N24 & N51 & N251 & N120; 
assign N312 = N70 | N49; 
assign N313 = N60 | N63 | N116 | N172 | N189 | N191 | N258 | N267; 
assign N314 = N104 | N238 | N290 | N86; 
assign N315 = N64 | N143 | N179 | N199 | N223 | N236 | N262 | N265; 
assign N316 = N106 & N147 & N148 & N150 & N166 & N241 & N297 & N176 & N302; 
assign N317 = N22 & N33 & N83 & N88 & N169 & N279 & N303; 
assign N318 = N43 | N162 | N272 | N284; 
assign N319 = N249 | N268 | N305 | N286; 
assign N320 = N296 | N310; 
assign N321 = N110 | N149 | N155 | N207 | N255 | N264 | N306 | N307; 
assign N322 = N260 & N278 & N316; 
assign N323 = N142 | N237 | N246 | N289 | N294; 
assign N324 = N67 | N203 | N253 | N299 | N311; 
assign N325 = N62 | N208 | N239; 
assign N326 = N154 & N184 & N274; 
assign N327 = ~(N306); 
assign N328 = ~(N39); 
assign N329 = N59 | N195 | N285; 
assign N330 = N312 | N313; 
assign N331 = N263 | N301 | N308; 
assign N332 = N295 & N317 & N288; 
assign N333 = N9 | N151 | N248 | N257; 
assign N334 = N213 | N269; 
assign N335 = N105 & N164 & N181 & N266 & N275 & N304; 
assign N336 = N108 | N180 | N240 | N276; 
assign N337 = N7 | N144 | N160 | N243 | N254; 
assign N338 = N95 | N173 | N298; 
assign N339 = N35 | N152 | N287 | N314 | N315; 
assign N340 = N76 & N174 & N225; 
assign N341 = N89 & N227 & N247 & N309; 
assign N342 = N170 & N250 & N293; 
endmodule
