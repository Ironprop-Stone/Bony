module Depth_10_20_Nodes_200_400_S007 (N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N286, N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297, N298, N299, N300, N301, N302, N303, N304, N305, N306);

input N1; 
input N2; 
input N3; 
input N4; 
input N5; 
input N6; 
input N7; 
input N8; 
input N9; 
input N10; 
input N11; 
input N12; 
input N13; 

output N286; 
output N287; 
output N288; 
output N289; 
output N290; 
output N291; 
output N292; 
output N293; 
output N294; 
output N295; 
output N296; 
output N297; 
output N298; 
output N299; 
output N300; 
output N301; 
output N302; 
output N303; 
output N304; 
output N305; 
output N306; 

wire N14; 
wire N15; 
wire N16; 
wire N17; 
wire N18; 
wire N19; 
wire N20; 
wire N21; 
wire N22; 
wire N23; 
wire N24; 
wire N25; 
wire N26; 
wire N27; 
wire N28; 
wire N29; 
wire N30; 
wire N31; 
wire N32; 
wire N33; 
wire N34; 
wire N35; 
wire N36; 
wire N37; 
wire N38; 
wire N39; 
wire N40; 
wire N41; 
wire N42; 
wire N43; 
wire N44; 
wire N45; 
wire N46; 
wire N47; 
wire N48; 
wire N49; 
wire N50; 
wire N51; 
wire N52; 
wire N53; 
wire N54; 
wire N55; 
wire N56; 
wire N57; 
wire N58; 
wire N59; 
wire N60; 
wire N61; 
wire N62; 
wire N63; 
wire N64; 
wire N65; 
wire N66; 
wire N67; 
wire N68; 
wire N69; 
wire N70; 
wire N71; 
wire N72; 
wire N73; 
wire N74; 
wire N75; 
wire N76; 
wire N77; 
wire N78; 
wire N79; 
wire N80; 
wire N81; 
wire N82; 
wire N83; 
wire N84; 
wire N85; 
wire N86; 
wire N87; 
wire N88; 
wire N89; 
wire N90; 
wire N91; 
wire N92; 
wire N93; 
wire N94; 
wire N95; 
wire N96; 
wire N97; 
wire N98; 
wire N99; 
wire N100; 
wire N101; 
wire N102; 
wire N103; 
wire N104; 
wire N105; 
wire N106; 
wire N107; 
wire N108; 
wire N109; 
wire N110; 
wire N111; 
wire N112; 
wire N113; 
wire N114; 
wire N115; 
wire N116; 
wire N117; 
wire N118; 
wire N119; 
wire N120; 
wire N121; 
wire N122; 
wire N123; 
wire N124; 
wire N125; 
wire N126; 
wire N127; 
wire N128; 
wire N129; 
wire N130; 
wire N131; 
wire N132; 
wire N133; 
wire N134; 
wire N135; 
wire N136; 
wire N137; 
wire N138; 
wire N139; 
wire N140; 
wire N141; 
wire N142; 
wire N143; 
wire N144; 
wire N145; 
wire N146; 
wire N147; 
wire N148; 
wire N149; 
wire N150; 
wire N151; 
wire N152; 
wire N153; 
wire N154; 
wire N155; 
wire N156; 
wire N157; 
wire N158; 
wire N159; 
wire N160; 
wire N161; 
wire N162; 
wire N163; 
wire N164; 
wire N165; 
wire N166; 
wire N167; 
wire N168; 
wire N169; 
wire N170; 
wire N171; 
wire N172; 
wire N173; 
wire N174; 
wire N175; 
wire N176; 
wire N177; 
wire N178; 
wire N179; 
wire N180; 
wire N181; 
wire N182; 
wire N183; 
wire N184; 
wire N185; 
wire N186; 
wire N187; 
wire N188; 
wire N189; 
wire N190; 
wire N191; 
wire N192; 
wire N193; 
wire N194; 
wire N195; 
wire N196; 
wire N197; 
wire N198; 
wire N199; 
wire N200; 
wire N201; 
wire N202; 
wire N203; 
wire N204; 
wire N205; 
wire N206; 
wire N207; 
wire N208; 
wire N209; 
wire N210; 
wire N211; 
wire N212; 
wire N213; 
wire N214; 
wire N215; 
wire N216; 
wire N217; 
wire N218; 
wire N219; 
wire N220; 
wire N221; 
wire N222; 
wire N223; 
wire N224; 
wire N225; 
wire N226; 
wire N227; 
wire N228; 
wire N229; 
wire N230; 
wire N231; 
wire N232; 
wire N233; 
wire N234; 
wire N235; 
wire N236; 
wire N237; 
wire N238; 
wire N239; 
wire N240; 
wire N241; 
wire N242; 
wire N243; 
wire N244; 
wire N245; 
wire N246; 
wire N247; 
wire N248; 
wire N249; 
wire N250; 
wire N251; 
wire N252; 
wire N253; 
wire N254; 
wire N255; 
wire N256; 
wire N257; 
wire N258; 
wire N259; 
wire N260; 
wire N261; 
wire N262; 
wire N263; 
wire N264; 
wire N265; 
wire N266; 
wire N267; 
wire N268; 
wire N269; 
wire N270; 
wire N271; 
wire N272; 
wire N273; 
wire N274; 
wire N275; 
wire N276; 
wire N277; 
wire N278; 
wire N279; 
wire N280; 
wire N281; 
wire N282; 
wire N283; 
wire N284; 
wire N285; 

assign N14 = ~(N8); 
assign N15 = ~(N7); 
assign N16 = ~(N10); 
assign N17 = ~(N9); 
assign N18 = N7 | N8; 
assign N19 = ~(N11); 
assign N20 = ~(N7); 
assign N21 = ~(N4); 
assign N22 = ~(N4); 
assign N23 = ~(N7); 
assign N24 = ~(N8); 
assign N25 = ~(N5); 
assign N26 = N5 | N25 | N4; 
assign N27 = N14 & N16; 
assign N28 = ~(N11); 
assign N29 = N19 | N24 | N6; 
assign N30 = ~(N18); 
assign N31 = ~(N27); 
assign N32 = ~(N4); 
assign N33 = ~(N9); 
assign N34 = N10 | N29; 
assign N35 = ~(N27); 
assign N36 = ~(N18); 
assign N37 = ~(N10); 
assign N38 = ~(N13); 
assign N39 = ~(N26); 
assign N40 = N17 & N7; 
assign N41 = N23 & N9; 
assign N42 = N22 & N26; 
assign N43 = N21 & N27 & N15; 
assign N44 = ~(N33); 
assign N45 = N11 & N30 & N37; 
assign N46 = N1 & N4 & N31; 
assign N47 = N8 & N9 & N20 & N41 & N30; 
assign N48 = N40 | N6; 
assign N49 = N28 & N40; 
assign N50 = ~(N26); 
assign N51 = N15 | N31 | N20; 
assign N52 = ~(N1); 
assign N53 = ~(N37); 
assign N54 = ~(N36); 
assign N55 = N13 & N29; 
assign N56 = ~(N3); 
assign N57 = N3 & N15; 
assign N58 = N32 | N36; 
assign N59 = N45 & N51; 
assign N60 = ~(N14); 
assign N61 = N43 & N44 & N47; 
assign N62 = N33 | N30; 
assign N63 = N52 | N27; 
assign N64 = ~(N57); 
assign N65 = N2 & N39 & N38; 
assign N66 = ~(N46); 
assign N67 = ~(N44); 
assign N68 = ~(N57); 
assign N69 = ~(N55); 
assign N70 = N12 & N11; 
assign N71 = ~(N44); 
assign N72 = N6 & N44; 
assign N73 = N29 | N34; 
assign N74 = ~(N53); 
assign N75 = ~(N6); 
assign N76 = ~(N20); 
assign N77 = ~(N23); 
assign N78 = ~(N32); 
assign N79 = N69 & N46; 
assign N80 = ~(N38); 
assign N81 = N67 | N29; 
assign N82 = N46 | N44; 
assign N83 = N38 & N28; 
assign N84 = ~(N48); 
assign N85 = ~(N51); 
assign N86 = N18 | N48 | N29; 
assign N87 = ~(N12); 
assign N88 = N26 & N32; 
assign N89 = N57 | N24; 
assign N90 = N82 | N3; 
assign N91 = N63 | N31; 
assign N92 = ~(N55); 
assign N93 = N36 & N60 & N61 & N33; 
assign N94 = N42 & N75 & N77 & N8; 
assign N95 = N68 | N43; 
assign N96 = N35 | N49 | N71 | N87 | N25; 
assign N97 = N34 & N70 & N45; 
assign N98 = ~(N44); 
assign N99 = N56 & N64 & N76 & N89 & N43; 
assign N100 = N47 | N74 | N93 | N96 | N58; 
assign N101 = ~(N53); 
assign N102 = N50 | N92 | N30; 
assign N103 = N53 | N58 | N79 | N3; 
assign N104 = N54 & N73 & N5; 
assign N105 = ~(N18); 
assign N106 = ~(N53); 
assign N107 = ~(N38); 
assign N108 = ~(N42); 
assign N109 = ~(N26); 
assign N110 = ~(N42); 
assign N111 = ~(N31); 
assign N112 = ~(N46); 
assign N113 = N55 | N65 | N43; 
assign N114 = ~(N43); 
assign N115 = ~(N10); 
assign N116 = N51 & N62 & N3; 
assign N117 = N81 & N40; 
assign N118 = ~(N21); 
assign N119 = ~(N19); 
assign N120 = ~(N53); 
assign N121 = ~(N56); 
assign N122 = N80 & N46; 
assign N123 = N91 & N100; 
assign N124 = ~(N35); 
assign N125 = ~(N59); 
assign N126 = ~(N20); 
assign N127 = ~(N90); 
assign N128 = ~(N15); 
assign N129 = ~(N27); 
assign N130 = ~(N24); 
assign N131 = ~(N23); 
assign N132 = ~(N45); 
assign N133 = ~(N69); 
assign N134 = ~(N55); 
assign N135 = ~(N22); 
assign N136 = ~(N22); 
assign N137 = ~(N50); 
assign N138 = ~(N84); 
assign N139 = ~(N45); 
assign N140 = N109 & N45; 
assign N141 = ~(N47); 
assign N142 = ~(N34); 
assign N143 = ~(N15); 
assign N144 = ~(N89); 
assign N145 = ~(N38); 
assign N146 = ~(N86); 
assign N147 = ~(N50); 
assign N148 = ~(N28); 
assign N149 = N115 | N55; 
assign N150 = ~(N28); 
assign N151 = N66 | N25; 
assign N152 = N106 & N54; 
assign N153 = ~(N28); 
assign N154 = ~(N1); 
assign N155 = ~(N101); 
assign N156 = N102 & N21; 
assign N157 = ~(N18); 
assign N158 = ~(N13); 
assign N159 = ~(N47); 
assign N160 = ~(N30); 
assign N161 = ~(N21); 
assign N162 = ~(N42); 
assign N163 = ~(N26); 
assign N164 = ~(N93); 
assign N165 = ~(N39); 
assign N166 = ~(N30); 
assign N167 = ~(N117); 
assign N168 = ~(N17); 
assign N169 = ~(N40); 
assign N170 = ~(N112); 
assign N171 = ~(N41); 
assign N172 = ~(N112); 
assign N173 = ~(N40); 
assign N174 = ~(N21); 
assign N175 = ~(N108); 
assign N176 = ~(N107); 
assign N177 = ~(N108); 
assign N178 = ~(N54); 
assign N179 = ~(N100); 
assign N180 = ~(N39); 
assign N181 = ~(N68); 
assign N182 = ~(N114); 
assign N183 = ~(N55); 
assign N184 = ~(N4); 
assign N185 = ~(N13); 
assign N186 = ~(N24); 
assign N187 = ~(N10); 
assign N188 = ~(N93); 
assign N189 = N118 & N1; 
assign N190 = ~(N85); 
assign N191 = ~(N106); 
assign N192 = N85 & N90; 
assign N193 = ~(N14); 
assign N194 = ~(N40); 
assign N195 = ~(N19); 
assign N196 = ~(N19); 
assign N197 = ~(N5); 
assign N198 = N83 & N49; 
assign N199 = N72 | N10; 
assign N200 = ~(N42); 
assign N201 = ~(N22); 
assign N202 = ~(N33); 
assign N203 = ~(N39); 
assign N204 = N111 & N158 & N194 & N42; 
assign N205 = ~(N94); 
assign N206 = N104 & N120 & N138 & N149; 
assign N207 = N183 | N184 | N47; 
assign N208 = N95 | N119 | N123 | N167 | N196 | N39; 
assign N209 = ~(N88); 
assign N210 = N121 & N201; 
assign N211 = N78 | N105 | N141 | N166; 
assign N212 = N84 | N99; 
assign N213 = N126 | N185; 
assign N214 = N162 | N51; 
assign N215 = ~(N47); 
assign N216 = ~(N97); 
assign N217 = N188 | N36; 
assign N218 = N101 & N207 & N212 & N215 & N19; 
assign N219 = N134 | N146 | N20; 
assign N220 = N156 | N164; 
assign N221 = N155 & N174 & N192 & N54; 
assign N222 = ~(N128); 
assign N223 = ~(N94); 
assign N224 = N129 & N172 & N32; 
assign N225 = ~(N98); 
assign N226 = N137 | N143 | N211 | N51; 
assign N227 = N168 | N31; 
assign N228 = ~(N176); 
assign N229 = ~(N84); 
assign N230 = N117 | N151; 
assign N231 = ~(N124); 
assign N232 = ~(N139); 
assign N233 = N110 & N58; 
assign N234 = ~(N175); 
assign N235 = N186 & N210 & N52; 
assign N236 = ~(N133); 
assign N237 = N144 & N161 & N163 & N204 & N220 & N236; 
assign N238 = N169 & N179 & N199 & N218 & N235; 
assign N239 = N127 & N130 & N178 & N191 & N206 & N221; 
assign N240 = N152 & N187 & N233 & N39; 
assign N241 = N160 & N195 & N213 & N231 & N24; 
assign N242 = N125 & N147 & N171 & N222 & N226 & N49; 
assign N243 = N132 & N209 & N36; 
assign N244 = ~(N103); 
assign N245 = ~(N205); 
assign N246 = N128 | N22; 
assign N247 = ~(N49); 
assign N248 = ~(N58); 
assign N249 = N170 | N193; 
assign N250 = ~(N116); 
assign N251 = ~(N165); 
assign N252 = ~(N23); 
assign N253 = N216 & N6; 
assign N254 = ~(N36); 
assign N255 = N148 | N150; 
assign N256 = ~(N17); 
assign N257 = ~(N49); 
assign N258 = ~(N215); 
assign N259 = ~(N202); 
assign N260 = ~(N81); 
assign N261 = ~(N1); 
assign N262 = ~(N160); 
assign N263 = ~(N140); 
assign N264 = ~(N208); 
assign N265 = ~(N35); 
assign N266 = ~(N14); 
assign N267 = ~(N131); 
assign N268 = ~(N119); 
assign N269 = N200 | N227 | N41; 
assign N270 = N157 & N177; 
assign N271 = ~(N33); 
assign N272 = ~(N23); 
assign N273 = N240 | N25; 
assign N274 = N182 | N54; 
assign N275 = N159 & N32; 
assign N276 = ~(N234); 
assign N277 = ~(N52); 
assign N278 = ~(N2); 
assign N279 = ~(N46); 
assign N280 = ~(N202); 
assign N281 = N135 & N230 & N52; 
assign N282 = ~(N48); 
assign N283 = ~(N181); 
assign N284 = ~(N11); 
assign N285 = ~(N23); 
assign N286 = N243 & N259 & N285; 
assign N287 = N107 & N153 & N203 & N251 & N263 & N283; 
assign N288 = N190 & N225 & N239 & N250 & N272; 
assign N289 = N142 | N246; 
assign N290 = N173 | N266; 
assign N291 = N122 | N282; 
assign N292 = N113 & N175 & N241 & N277 & N284; 
assign N293 = N229 | N242 | N268; 
assign N294 = N116 & N232 & N257 & N265 & N278; 
assign N295 = N228 | N270 | N273; 
assign N296 = ~(N279); 
assign N297 = N198 | N248 | N252 | N260 | N274; 
assign N298 = N136 & N269 & N276; 
assign N299 = N244 | N247 | N275; 
assign N300 = N189 | N253 | N258 | N271; 
assign N301 = N154 | N219 | N238 | N256; 
assign N302 = N205 & N217 & N249 & N264 & N280; 
assign N303 = N180 & N214 & N224 & N254 & N262; 
assign N304 = N237 & N245 & N255; 
assign N305 = N197 & N261 & N267; 
assign N306 = N145 & N223 & N281; 
endmodule
