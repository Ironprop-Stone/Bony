module Depth_10_20_Nodes_200_400_S003 (N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N322, N323, N324, N325, N326, N327, N328, N329, N330, N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341, N342, N343, N344);

input N1; 
input N2; 
input N3; 
input N4; 
input N5; 
input N6; 
input N7; 
input N8; 
input N9; 
input N10; 
input N11; 
input N12; 
input N13; 
input N14; 
input N15; 
input N16; 

output N322; 
output N323; 
output N324; 
output N325; 
output N326; 
output N327; 
output N328; 
output N329; 
output N330; 
output N331; 
output N332; 
output N333; 
output N334; 
output N335; 
output N336; 
output N337; 
output N338; 
output N339; 
output N340; 
output N341; 
output N342; 
output N343; 
output N344; 

wire N17; 
wire N18; 
wire N19; 
wire N20; 
wire N21; 
wire N22; 
wire N23; 
wire N24; 
wire N25; 
wire N26; 
wire N27; 
wire N28; 
wire N29; 
wire N30; 
wire N31; 
wire N32; 
wire N33; 
wire N34; 
wire N35; 
wire N36; 
wire N37; 
wire N38; 
wire N39; 
wire N40; 
wire N41; 
wire N42; 
wire N43; 
wire N44; 
wire N45; 
wire N46; 
wire N47; 
wire N48; 
wire N49; 
wire N50; 
wire N51; 
wire N52; 
wire N53; 
wire N54; 
wire N55; 
wire N56; 
wire N57; 
wire N58; 
wire N59; 
wire N60; 
wire N61; 
wire N62; 
wire N63; 
wire N64; 
wire N65; 
wire N66; 
wire N67; 
wire N68; 
wire N69; 
wire N70; 
wire N71; 
wire N72; 
wire N73; 
wire N74; 
wire N75; 
wire N76; 
wire N77; 
wire N78; 
wire N79; 
wire N80; 
wire N81; 
wire N82; 
wire N83; 
wire N84; 
wire N85; 
wire N86; 
wire N87; 
wire N88; 
wire N89; 
wire N90; 
wire N91; 
wire N92; 
wire N93; 
wire N94; 
wire N95; 
wire N96; 
wire N97; 
wire N98; 
wire N99; 
wire N100; 
wire N101; 
wire N102; 
wire N103; 
wire N104; 
wire N105; 
wire N106; 
wire N107; 
wire N108; 
wire N109; 
wire N110; 
wire N111; 
wire N112; 
wire N113; 
wire N114; 
wire N115; 
wire N116; 
wire N117; 
wire N118; 
wire N119; 
wire N120; 
wire N121; 
wire N122; 
wire N123; 
wire N124; 
wire N125; 
wire N126; 
wire N127; 
wire N128; 
wire N129; 
wire N130; 
wire N131; 
wire N132; 
wire N133; 
wire N134; 
wire N135; 
wire N136; 
wire N137; 
wire N138; 
wire N139; 
wire N140; 
wire N141; 
wire N142; 
wire N143; 
wire N144; 
wire N145; 
wire N146; 
wire N147; 
wire N148; 
wire N149; 
wire N150; 
wire N151; 
wire N152; 
wire N153; 
wire N154; 
wire N155; 
wire N156; 
wire N157; 
wire N158; 
wire N159; 
wire N160; 
wire N161; 
wire N162; 
wire N163; 
wire N164; 
wire N165; 
wire N166; 
wire N167; 
wire N168; 
wire N169; 
wire N170; 
wire N171; 
wire N172; 
wire N173; 
wire N174; 
wire N175; 
wire N176; 
wire N177; 
wire N178; 
wire N179; 
wire N180; 
wire N181; 
wire N182; 
wire N183; 
wire N184; 
wire N185; 
wire N186; 
wire N187; 
wire N188; 
wire N189; 
wire N190; 
wire N191; 
wire N192; 
wire N193; 
wire N194; 
wire N195; 
wire N196; 
wire N197; 
wire N198; 
wire N199; 
wire N200; 
wire N201; 
wire N202; 
wire N203; 
wire N204; 
wire N205; 
wire N206; 
wire N207; 
wire N208; 
wire N209; 
wire N210; 
wire N211; 
wire N212; 
wire N213; 
wire N214; 
wire N215; 
wire N216; 
wire N217; 
wire N218; 
wire N219; 
wire N220; 
wire N221; 
wire N222; 
wire N223; 
wire N224; 
wire N225; 
wire N226; 
wire N227; 
wire N228; 
wire N229; 
wire N230; 
wire N231; 
wire N232; 
wire N233; 
wire N234; 
wire N235; 
wire N236; 
wire N237; 
wire N238; 
wire N239; 
wire N240; 
wire N241; 
wire N242; 
wire N243; 
wire N244; 
wire N245; 
wire N246; 
wire N247; 
wire N248; 
wire N249; 
wire N250; 
wire N251; 
wire N252; 
wire N253; 
wire N254; 
wire N255; 
wire N256; 
wire N257; 
wire N258; 
wire N259; 
wire N260; 
wire N261; 
wire N262; 
wire N263; 
wire N264; 
wire N265; 
wire N266; 
wire N267; 
wire N268; 
wire N269; 
wire N270; 
wire N271; 
wire N272; 
wire N273; 
wire N274; 
wire N275; 
wire N276; 
wire N277; 
wire N278; 
wire N279; 
wire N280; 
wire N281; 
wire N282; 
wire N283; 
wire N284; 
wire N285; 
wire N286; 
wire N287; 
wire N288; 
wire N289; 
wire N290; 
wire N291; 
wire N292; 
wire N293; 
wire N294; 
wire N295; 
wire N296; 
wire N297; 
wire N298; 
wire N299; 
wire N300; 
wire N301; 
wire N302; 
wire N303; 
wire N304; 
wire N305; 
wire N306; 
wire N307; 
wire N308; 
wire N309; 
wire N310; 
wire N311; 
wire N312; 
wire N313; 
wire N314; 
wire N315; 
wire N316; 
wire N317; 
wire N318; 
wire N319; 
wire N320; 
wire N321; 

assign N17 = ~(N8); 
assign N18 = ~(N6); 
assign N19 = ~(N6); 
assign N20 = N6 | N1; 
assign N21 = ~(N10); 
assign N22 = ~(N10); 
assign N23 = ~(N14); 
assign N24 = ~(N15); 
assign N25 = ~(N6); 
assign N26 = ~(N5); 
assign N27 = ~(N9); 
assign N28 = N8 & N7; 
assign N29 = ~(N1); 
assign N30 = ~(N2); 
assign N31 = ~(N11); 
assign N32 = ~(N13); 
assign N33 = ~(N4); 
assign N34 = ~(N8); 
assign N35 = ~(N6); 
assign N36 = ~(N3); 
assign N37 = ~(N14); 
assign N38 = ~(N13); 
assign N39 = ~(N5); 
assign N40 = ~(N16); 
assign N41 = N15 & N10; 
assign N42 = ~(N5); 
assign N43 = ~(N8); 
assign N44 = ~(N1); 
assign N45 = ~(N12); 
assign N46 = ~(N15); 
assign N47 = ~(N9); 
assign N48 = ~(N13); 
assign N49 = ~(N12); 
assign N50 = ~(N15); 
assign N51 = ~(N1); 
assign N52 = ~(N5); 
assign N53 = ~(N13); 
assign N54 = ~(N4); 
assign N55 = ~(N7); 
assign N56 = ~(N8); 
assign N57 = N9 | N16; 
assign N58 = ~(N16); 
assign N59 = ~(N2); 
assign N60 = ~(N21); 
assign N61 = N35 & N44 & N2; 
assign N62 = ~(N12); 
assign N63 = ~(N16); 
assign N64 = ~(N14); 
assign N65 = N26 | N56; 
assign N66 = ~(N37); 
assign N67 = ~(N2); 
assign N68 = N46 & N31; 
assign N69 = N32 & N30; 
assign N70 = N30 & N3; 
assign N71 = ~(N12); 
assign N72 = N22 | N43; 
assign N73 = ~(N32); 
assign N74 = ~(N40); 
assign N75 = N61 | N34; 
assign N76 = ~(N15); 
assign N77 = ~(N66); 
assign N78 = ~(N9); 
assign N79 = ~(N43); 
assign N80 = ~(N4); 
assign N81 = ~(N64); 
assign N82 = ~(N4); 
assign N83 = N60 & N69 & N30; 
assign N84 = ~(N63); 
assign N85 = ~(N27); 
assign N86 = N67 & N61; 
assign N87 = N4 & N48; 
assign N88 = ~(N70); 
assign N89 = N42 & N49; 
assign N90 = N53 & N55 & N14; 
assign N91 = ~(N35); 
assign N92 = N50 | N88; 
assign N93 = N49 | N40; 
assign N94 = ~(N66); 
assign N95 = ~(N65); 
assign N96 = ~(N12); 
assign N97 = N10 | N39 | N48 | N44; 
assign N98 = N23 | N59 | N87; 
assign N99 = N7 & N51 & N76 & N11; 
assign N100 = ~(N83); 
assign N101 = ~(N63); 
assign N102 = N13 | N10; 
assign N103 = ~(N70); 
assign N104 = ~(N68); 
assign N105 = N68 | N21; 
assign N106 = N45 & N70; 
assign N107 = ~(N55); 
assign N108 = N21 & N28 & N33 & N36 & N3; 
assign N109 = N20 & N89 & N99; 
assign N110 = N5 & N11 & N47 & N63 & N71 & N102 & N86; 
assign N111 = N2 | N38 | N77 | N93; 
assign N112 = N1 & N29; 
assign N113 = ~(N95); 
assign N114 = N14 | N84 | N105; 
assign N115 = N18 | N19 | N57 | N76; 
assign N116 = ~(N65); 
assign N117 = ~(N75); 
assign N118 = N31 | N92 | N106; 
assign N119 = N74 & N30; 
assign N120 = N75 & N89; 
assign N121 = N17 & N83 & N65; 
assign N122 = N3 | N61; 
assign N123 = ~(N5); 
assign N124 = ~(N66); 
assign N125 = N91 & N64; 
assign N126 = ~(N108); 
assign N127 = N16 | N41 | N88 | N101 | N106 | N61; 
assign N128 = N82 | N101; 
assign N129 = N96 | N55; 
assign N130 = N111 & N103; 
assign N131 = ~(N108); 
assign N132 = N34 | N97 | N112; 
assign N133 = N66 | N70 | N25; 
assign N134 = N25 | N64; 
assign N135 = N52 & N90 & N103 & N112; 
assign N136 = N56 & N58 & N103; 
assign N137 = ~(N88); 
assign N138 = ~(N104); 
assign N139 = N24 & N113 & N98; 
assign N140 = ~(N93); 
assign N141 = N62 & N85; 
assign N142 = ~(N123); 
assign N143 = N119 | N111; 
assign N144 = ~(N107); 
assign N145 = N65 | N110; 
assign N146 = ~(N95); 
assign N147 = N40 & N54 & N98 & N96; 
assign N148 = N93 & N68; 
assign N149 = ~(N77); 
assign N150 = ~(N91); 
assign N151 = N124 & N27; 
assign N152 = ~(N109); 
assign N153 = N117 & N91; 
assign N154 = ~(N16); 
assign N155 = ~(N57); 
assign N156 = ~(N105); 
assign N157 = ~(N84); 
assign N158 = ~(N82); 
assign N159 = ~(N21); 
assign N160 = ~(N90); 
assign N161 = ~(N69); 
assign N162 = N79 & N80 & N94 & N19; 
assign N163 = N85 | N107; 
assign N164 = ~(N98); 
assign N165 = ~(N65); 
assign N166 = N73 & N105; 
assign N167 = ~(N92); 
assign N168 = N72 & N108; 
assign N169 = ~(N116); 
assign N170 = ~(N107); 
assign N171 = ~(N68); 
assign N172 = N81 | N70; 
assign N173 = ~(N97); 
assign N174 = N116 | N98; 
assign N175 = ~(N108); 
assign N176 = N129 | N135 | N91; 
assign N177 = ~(N36); 
assign N178 = ~(N23); 
assign N179 = N115 | N37; 
assign N180 = ~(N81); 
assign N181 = ~(N69); 
assign N182 = N78 & N104; 
assign N183 = ~(N108); 
assign N184 = ~(N45); 
assign N185 = ~(N7); 
assign N186 = ~(N103); 
assign N187 = ~(N93); 
assign N188 = ~(N69); 
assign N189 = N64 | N109; 
assign N190 = ~(N83); 
assign N191 = ~(N109); 
assign N192 = ~(N80); 
assign N193 = N187 & N33; 
assign N194 = N87 | N95; 
assign N195 = ~(N159); 
assign N196 = N86 | N109; 
assign N197 = ~(N108); 
assign N198 = N168 | N186 | N71; 
assign N199 = N139 | N63; 
assign N200 = N120 | N68; 
assign N201 = N141 & N147 & N169 & N189 & N82; 
assign N202 = N130 | N2; 
assign N203 = N95 | N170 | N109; 
assign N204 = N164 & N44; 
assign N205 = N100 & N121 & N150 & N158 & N165 & N179 & N41; 
assign N206 = N185 | N61; 
assign N207 = N131 & N161 & N44; 
assign N208 = N112 & N114 & N125 & N71; 
assign N209 = N167 & N47; 
assign N210 = ~(N40); 
assign N211 = N99 & N153 & N159 & N194 & N77; 
assign N212 = N151 & N82; 
assign N213 = N172 & N104; 
assign N214 = N132 & N191 & N101; 
assign N215 = ~(N104); 
assign N216 = ~(N73); 
assign N217 = N178 | N90; 
assign N218 = N133 & N137 & N144 & N197 & N55; 
assign N219 = N110 | N163 | N69; 
assign N220 = N181 & N11; 
assign N221 = ~(N44); 
assign N222 = ~(N9); 
assign N223 = N107 & N88; 
assign N224 = N122 | N127 | N34; 
assign N225 = N140 | N107; 
assign N226 = ~(N85); 
assign N227 = ~(N91); 
assign N228 = ~(N148); 
assign N229 = N123 | N173 | N184 | N211 | N224 | N63; 
assign N230 = N126 & N209; 
assign N231 = N142 & N155 & N106; 
assign N232 = N118 | N75; 
assign N233 = N160 & N218 & N223 & N73; 
assign N234 = N149 | N177 | N86; 
assign N235 = N174 & N180 & N195 & N200 & N216 & N27; 
assign N236 = N128 & N154 & N156 & N43; 
assign N237 = N176 | N204 | N208; 
assign N238 = N152 | N89; 
assign N239 = N134 | N138 | N143 | N145 | N220 | N231 | N77; 
assign N240 = N136 & N175 & N104; 
assign N241 = N146 | N171 | N206 | N112; 
assign N242 = N190 | N199 | N80; 
assign N243 = ~(N111); 
assign N244 = ~(N95); 
assign N245 = ~(N111); 
assign N246 = ~(N140); 
assign N247 = N215 & N228 & N60; 
assign N248 = N157 & N192 & N37; 
assign N249 = ~(N49); 
assign N250 = ~(N237); 
assign N251 = ~(N72); 
assign N252 = ~(N36); 
assign N253 = N205 | N110; 
assign N254 = ~(N40); 
assign N255 = ~(N28); 
assign N256 = ~(N242); 
assign N257 = ~(N74); 
assign N258 = ~(N106); 
assign N259 = ~(N87); 
assign N260 = ~(N42); 
assign N261 = ~(N215); 
assign N262 = ~(N112); 
assign N263 = ~(N222); 
assign N264 = ~(N241); 
assign N265 = N162 & N94; 
assign N266 = ~(N182); 
assign N267 = ~(N210); 
assign N268 = N166 & N201 & N87; 
assign N269 = N233 & N32; 
assign N270 = ~(N133); 
assign N271 = ~(N221); 
assign N272 = ~(N183); 
assign N273 = ~(N79); 
assign N274 = ~(N80); 
assign N275 = N188 & N106; 
assign N276 = N212 & N219 & N240 & N253 & N58; 
assign N277 = N251 & N263; 
assign N278 = N198 | N207 | N225 | N232 | N247 | N87; 
assign N279 = N193 | N246 | N264 | N86; 
assign N280 = N196 | N202 | N226 | N270 | N106; 
assign N281 = N262 & N92; 
assign N282 = ~(N97); 
assign N283 = ~(N33); 
assign N284 = N229 & N111; 
assign N285 = N255 & N17; 
assign N286 = N239 & N71; 
assign N287 = ~(N68); 
assign N288 = N258 | N7; 
assign N289 = N222 & N227 & N254 & N275; 
assign N290 = N249 | N257 | N71; 
assign N291 = N203 | N280 | N105; 
assign N292 = ~(N3); 
assign N293 = ~(N107); 
assign N294 = ~(N58); 
assign N295 = ~(N19); 
assign N296 = ~(N131); 
assign N297 = ~(N47); 
assign N298 = ~(N273); 
assign N299 = N279 | N81; 
assign N300 = ~(N224); 
assign N301 = ~(N235); 
assign N302 = ~(N31); 
assign N303 = ~(N213); 
assign N304 = ~(N256); 
assign N305 = ~(N103); 
assign N306 = N271 | N283 | N293; 
assign N307 = N236 & N245 & N261 & N299 & N11; 
assign N308 = N298 & N302 & N70; 
assign N309 = N265 & N294; 
assign N310 = N248 & N260 & N295; 
assign N311 = N284 & N289 & N90; 
assign N312 = N217 | N241; 
assign N313 = N274 | N277 | N285; 
assign N314 = N243 & N250 & N296 & N81; 
assign N315 = ~(N137); 
assign N316 = N214 | N244 | N259 | N266 | N269 | N282; 
assign N317 = N230 | N234 | N281 | N110; 
assign N318 = ~(N93); 
assign N319 = N287 & N300 & N20; 
assign N320 = ~(N80); 
assign N321 = ~(N101); 
assign N322 = ~(N54); 
assign N323 = N268 & N307 & N311; 
assign N324 = ~(N235); 
assign N325 = ~(N312); 
assign N326 = ~(N321); 
assign N327 = ~(N189); 
assign N328 = ~(N278); 
assign N329 = ~(N231); 
assign N330 = ~(N316); 
assign N331 = N303 | N308 | N314; 
assign N332 = N301 & N304 & N315; 
assign N333 = ~(N317); 
assign N334 = ~(N286); 
assign N335 = N292 & N306 & N318; 
assign N336 = N267 & N290 & N313; 
assign N337 = N238 & N305; 
assign N338 = ~(N278); 
assign N339 = N288 | N291 | N297; 
assign N340 = ~(N118); 
assign N341 = ~(N237); 
assign N342 = ~(N207); 
assign N343 = N252 & N310 & N319 & N320; 
assign N344 = N272 & N276 & N309; 
endmodule
