module test_00 (N1, N2, N3, N4, N34, N35, N36, N37, N38, N39, N40);

input N1; 
input N2; 
input N3; 
input N4; 

output N34; 
output N35; 
output N36; 
output N37; 
output N38; 
output N39; 
output N40; 

wire N5; 
wire N6; 
wire N7; 
wire N8; 
wire N9; 
wire N10; 
wire N11; 
wire N12; 
wire N13; 
wire N14; 
wire N15; 
wire N16; 
wire N17; 
wire N18; 
wire N19; 
wire N20; 
wire N21; 
wire N22; 
wire N23; 
wire N24; 
wire N25; 
wire N26; 
wire N27; 
wire N28; 
wire N29; 
wire N30; 
wire N31; 
wire N32; 
wire N33; 

assign N5 = N3 | N1; 
assign N6 = ~(N2); 
assign N7 = ~(N3); 
assign N8 = ~(N3); 
assign N9 = ~(N4); 
assign N10 = ~(N2); 
assign N11 = N2 | N5 | N6; 
assign N12 = ~(N8); 
assign N13 = ~(N8); 
assign N14 = ~(N5); 
assign N15 = ~(N1); 
assign N16 = N7 | N8 | N2; 
assign N17 = ~(N4); 
assign N18 = N6 | N12 | N4; 
assign N19 = N1 | N10; 
assign N20 = ~(N3); 
assign N21 = ~(N2); 
assign N22 = N15 | N17; 
assign N23 = N14 & N10 & N9 & N18 & N15 & N12 & N17 & N6 & N13; 
assign N24 = N10 & N16 & N5; 
assign N25 = ~(N12); 
assign N26 = ~(N15); 
assign N27 = N20 & N23 & N15; 
assign N28 = ~(N3); 
assign N29 = ~(N4); 
assign N30 = ~(N25); 
assign N31 = N13 | N24 | N29 | N23; 
assign N32 = N21 | N30; 
assign N33 = N25 & N28 & N30 & N4; 
assign N34 = ~(N18); 
assign N35 = N14 | N27 | N32; 
assign N36 = N22 | N31; 
assign N37 = N16 & N18 & N1 & N32 & N14 & N29 & N15 & N7 & N11; 
assign N38 = ~(N11); 
assign N39 = N9 & N19 & N26 & N33; 
assign N40 = ~(N17); 
endmodule
