module test_02 (N1, N2, N3, N4, N5, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42);

input N1; 
input N2; 
input N3; 
input N4; 
input N5; 

output N32; 
output N33; 
output N34; 
output N35; 
output N36; 
output N37; 
output N38; 
output N39; 
output N40; 
output N41; 
output N42; 

wire N6; 
wire N7; 
wire N8; 
wire N9; 
wire N10; 
wire N11; 
wire N12; 
wire N13; 
wire N14; 
wire N15; 
wire N16; 
wire N17; 
wire N18; 
wire N19; 
wire N20; 
wire N21; 
wire N22; 
wire N23; 
wire N24; 
wire N25; 
wire N26; 
wire N27; 
wire N28; 
wire N29; 
wire N30; 
wire N31; 

assign N6 = ~(N1); 
assign N7 = ~(N2); 
assign N8 = ~(N2); 
assign N9 = ~(N3); 
assign N10 = ~(N1); 
assign N11 = ~(N3); 
assign N12 = ~(N3); 
assign N13 = ~(N2); 
assign N14 = ~(N2); 
assign N15 = ~(N4); 
assign N16 = ~(N3); 
assign N17 = N10 | N5; 
assign N18 = N14 & N7; 
assign N19 = N12 | N13; 
assign N20 = ~(N5); 
assign N21 = N13 & N1; 
assign N22 = ~(N10); 
assign N23 = N20 | N9; 
assign N24 = ~(N1); 
assign N25 = N1 | N12; 
assign N26 = ~(N19); 
assign N27 = N5 | N18 | N4 | N1 | N2 | N3 | N12 | N17 | N16; 
assign N28 = N3 & N8 & N19 & N27; 
assign N29 = N11 & N15 & N21 & N23 & N26; 
assign N30 = N4 & N9 & N24; 
assign N31 = N16 & N25 & N21; 
assign N32 = N21 & N22 & N9 & N19 & N25 & N4 & N10 & N28 & N8; 
assign N33 = N29 | N31; 
assign N34 = N21 & N30 & N14 & N22 & N4 & N31 & N29 & N25 & N18; 
assign N35 = N31 & N29 & N6 & N30 & N27 & N16 & N10 & N17 & N14; 
assign N36 = ~(N17); 
assign N37 = ~(N18); 
assign N38 = N5 | N7 | N28 | N30; 
assign N39 = ~(N22); 
assign N40 = ~(N2); 
assign N41 = ~(N6); 
assign N42 = N4 & N30 & N23 & N7 & N28 & N29 & N17 & N31 & N26; 
endmodule
