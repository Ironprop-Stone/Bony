module Depth_10_20_Nodes_200_400_S001 (N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N444, N445, N446, N447, N448, N449, N450, N451, N452, N453, N454, N455, N456, N457, N458, N459, N460, N461, N462, N463, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473, N474, N475, N476, N477, N478, N479, N480, N481);

input N1; 
input N2; 
input N3; 
input N4; 
input N5; 
input N6; 
input N7; 
input N8; 
input N9; 
input N10; 
input N11; 
input N12; 
input N13; 
input N14; 
input N15; 

output N444; 
output N445; 
output N446; 
output N447; 
output N448; 
output N449; 
output N450; 
output N451; 
output N452; 
output N453; 
output N454; 
output N455; 
output N456; 
output N457; 
output N458; 
output N459; 
output N460; 
output N461; 
output N462; 
output N463; 
output N464; 
output N465; 
output N466; 
output N467; 
output N468; 
output N469; 
output N470; 
output N471; 
output N472; 
output N473; 
output N474; 
output N475; 
output N476; 
output N477; 
output N478; 
output N479; 
output N480; 
output N481; 

wire N16; 
wire N17; 
wire N18; 
wire N19; 
wire N20; 
wire N21; 
wire N22; 
wire N23; 
wire N24; 
wire N25; 
wire N26; 
wire N27; 
wire N28; 
wire N29; 
wire N30; 
wire N31; 
wire N32; 
wire N33; 
wire N34; 
wire N35; 
wire N36; 
wire N37; 
wire N38; 
wire N39; 
wire N40; 
wire N41; 
wire N42; 
wire N43; 
wire N44; 
wire N45; 
wire N46; 
wire N47; 
wire N48; 
wire N49; 
wire N50; 
wire N51; 
wire N52; 
wire N53; 
wire N54; 
wire N55; 
wire N56; 
wire N57; 
wire N58; 
wire N59; 
wire N60; 
wire N61; 
wire N62; 
wire N63; 
wire N64; 
wire N65; 
wire N66; 
wire N67; 
wire N68; 
wire N69; 
wire N70; 
wire N71; 
wire N72; 
wire N73; 
wire N74; 
wire N75; 
wire N76; 
wire N77; 
wire N78; 
wire N79; 
wire N80; 
wire N81; 
wire N82; 
wire N83; 
wire N84; 
wire N85; 
wire N86; 
wire N87; 
wire N88; 
wire N89; 
wire N90; 
wire N91; 
wire N92; 
wire N93; 
wire N94; 
wire N95; 
wire N96; 
wire N97; 
wire N98; 
wire N99; 
wire N100; 
wire N101; 
wire N102; 
wire N103; 
wire N104; 
wire N105; 
wire N106; 
wire N107; 
wire N108; 
wire N109; 
wire N110; 
wire N111; 
wire N112; 
wire N113; 
wire N114; 
wire N115; 
wire N116; 
wire N117; 
wire N118; 
wire N119; 
wire N120; 
wire N121; 
wire N122; 
wire N123; 
wire N124; 
wire N125; 
wire N126; 
wire N127; 
wire N128; 
wire N129; 
wire N130; 
wire N131; 
wire N132; 
wire N133; 
wire N134; 
wire N135; 
wire N136; 
wire N137; 
wire N138; 
wire N139; 
wire N140; 
wire N141; 
wire N142; 
wire N143; 
wire N144; 
wire N145; 
wire N146; 
wire N147; 
wire N148; 
wire N149; 
wire N150; 
wire N151; 
wire N152; 
wire N153; 
wire N154; 
wire N155; 
wire N156; 
wire N157; 
wire N158; 
wire N159; 
wire N160; 
wire N161; 
wire N162; 
wire N163; 
wire N164; 
wire N165; 
wire N166; 
wire N167; 
wire N168; 
wire N169; 
wire N170; 
wire N171; 
wire N172; 
wire N173; 
wire N174; 
wire N175; 
wire N176; 
wire N177; 
wire N178; 
wire N179; 
wire N180; 
wire N181; 
wire N182; 
wire N183; 
wire N184; 
wire N185; 
wire N186; 
wire N187; 
wire N188; 
wire N189; 
wire N190; 
wire N191; 
wire N192; 
wire N193; 
wire N194; 
wire N195; 
wire N196; 
wire N197; 
wire N198; 
wire N199; 
wire N200; 
wire N201; 
wire N202; 
wire N203; 
wire N204; 
wire N205; 
wire N206; 
wire N207; 
wire N208; 
wire N209; 
wire N210; 
wire N211; 
wire N212; 
wire N213; 
wire N214; 
wire N215; 
wire N216; 
wire N217; 
wire N218; 
wire N219; 
wire N220; 
wire N221; 
wire N222; 
wire N223; 
wire N224; 
wire N225; 
wire N226; 
wire N227; 
wire N228; 
wire N229; 
wire N230; 
wire N231; 
wire N232; 
wire N233; 
wire N234; 
wire N235; 
wire N236; 
wire N237; 
wire N238; 
wire N239; 
wire N240; 
wire N241; 
wire N242; 
wire N243; 
wire N244; 
wire N245; 
wire N246; 
wire N247; 
wire N248; 
wire N249; 
wire N250; 
wire N251; 
wire N252; 
wire N253; 
wire N254; 
wire N255; 
wire N256; 
wire N257; 
wire N258; 
wire N259; 
wire N260; 
wire N261; 
wire N262; 
wire N263; 
wire N264; 
wire N265; 
wire N266; 
wire N267; 
wire N268; 
wire N269; 
wire N270; 
wire N271; 
wire N272; 
wire N273; 
wire N274; 
wire N275; 
wire N276; 
wire N277; 
wire N278; 
wire N279; 
wire N280; 
wire N281; 
wire N282; 
wire N283; 
wire N284; 
wire N285; 
wire N286; 
wire N287; 
wire N288; 
wire N289; 
wire N290; 
wire N291; 
wire N292; 
wire N293; 
wire N294; 
wire N295; 
wire N296; 
wire N297; 
wire N298; 
wire N299; 
wire N300; 
wire N301; 
wire N302; 
wire N303; 
wire N304; 
wire N305; 
wire N306; 
wire N307; 
wire N308; 
wire N309; 
wire N310; 
wire N311; 
wire N312; 
wire N313; 
wire N314; 
wire N315; 
wire N316; 
wire N317; 
wire N318; 
wire N319; 
wire N320; 
wire N321; 
wire N322; 
wire N323; 
wire N324; 
wire N325; 
wire N326; 
wire N327; 
wire N328; 
wire N329; 
wire N330; 
wire N331; 
wire N332; 
wire N333; 
wire N334; 
wire N335; 
wire N336; 
wire N337; 
wire N338; 
wire N339; 
wire N340; 
wire N341; 
wire N342; 
wire N343; 
wire N344; 
wire N345; 
wire N346; 
wire N347; 
wire N348; 
wire N349; 
wire N350; 
wire N351; 
wire N352; 
wire N353; 
wire N354; 
wire N355; 
wire N356; 
wire N357; 
wire N358; 
wire N359; 
wire N360; 
wire N361; 
wire N362; 
wire N363; 
wire N364; 
wire N365; 
wire N366; 
wire N367; 
wire N368; 
wire N369; 
wire N370; 
wire N371; 
wire N372; 
wire N373; 
wire N374; 
wire N375; 
wire N376; 
wire N377; 
wire N378; 
wire N379; 
wire N380; 
wire N381; 
wire N382; 
wire N383; 
wire N384; 
wire N385; 
wire N386; 
wire N387; 
wire N388; 
wire N389; 
wire N390; 
wire N391; 
wire N392; 
wire N393; 
wire N394; 
wire N395; 
wire N396; 
wire N397; 
wire N398; 
wire N399; 
wire N400; 
wire N401; 
wire N402; 
wire N403; 
wire N404; 
wire N405; 
wire N406; 
wire N407; 
wire N408; 
wire N409; 
wire N410; 
wire N411; 
wire N412; 
wire N413; 
wire N414; 
wire N415; 
wire N416; 
wire N417; 
wire N418; 
wire N419; 
wire N420; 
wire N421; 
wire N422; 
wire N423; 
wire N424; 
wire N425; 
wire N426; 
wire N427; 
wire N428; 
wire N429; 
wire N430; 
wire N431; 
wire N432; 
wire N433; 
wire N434; 
wire N435; 
wire N436; 
wire N437; 
wire N438; 
wire N439; 
wire N440; 
wire N441; 
wire N442; 
wire N443; 

assign N16 = ~(N2); 
assign N17 = ~(N10); 
assign N18 = ~(N4); 
assign N19 = ~(N3); 
assign N20 = ~(N12); 
assign N21 = ~(N5); 
assign N22 = ~(N6); 
assign N23 = ~(N13); 
assign N24 = ~(N12); 
assign N25 = ~(N8); 
assign N26 = ~(N12); 
assign N27 = ~(N10); 
assign N28 = ~(N10); 
assign N29 = ~(N15); 
assign N30 = ~(N11); 
assign N31 = N5 & N11; 
assign N32 = ~(N10); 
assign N33 = ~(N5); 
assign N34 = ~(N5); 
assign N35 = ~(N7); 
assign N36 = ~(N12); 
assign N37 = ~(N6); 
assign N38 = ~(N14); 
assign N39 = ~(N9); 
assign N40 = ~(N15); 
assign N41 = ~(N39); 
assign N42 = ~(N29); 
assign N43 = ~(N5); 
assign N44 = ~(N19); 
assign N45 = ~(N21); 
assign N46 = ~(N18); 
assign N47 = ~(N13); 
assign N48 = ~(N29); 
assign N49 = ~(N27); 
assign N50 = ~(N27); 
assign N51 = ~(N26); 
assign N52 = ~(N31); 
assign N53 = ~(N37); 
assign N54 = ~(N18); 
assign N55 = ~(N19); 
assign N56 = ~(N9); 
assign N57 = ~(N20); 
assign N58 = ~(N3); 
assign N59 = ~(N15); 
assign N60 = ~(N15); 
assign N61 = ~(N24); 
assign N62 = ~(N7); 
assign N63 = ~(N29); 
assign N64 = ~(N14); 
assign N65 = ~(N3); 
assign N66 = N35 & N40; 
assign N67 = N37 & N31; 
assign N68 = ~(N14); 
assign N69 = ~(N1); 
assign N70 = ~(N4); 
assign N71 = ~(N23); 
assign N72 = N29 | N1; 
assign N73 = ~(N21); 
assign N74 = ~(N27); 
assign N75 = ~(N25); 
assign N76 = N3 | N24; 
assign N77 = ~(N21); 
assign N78 = ~(N37); 
assign N79 = N31 | N41; 
assign N80 = ~(N23); 
assign N81 = N57 | N16; 
assign N82 = ~(N8); 
assign N83 = N55 & N76; 
assign N84 = ~(N54); 
assign N85 = N45 | N56; 
assign N86 = N64 & N65; 
assign N87 = N71 | N59; 
assign N88 = N22 | N52; 
assign N89 = ~(N76); 
assign N90 = ~(N47); 
assign N91 = ~(N51); 
assign N92 = ~(N1); 
assign N93 = ~(N64); 
assign N94 = ~(N79); 
assign N95 = N63 | N74; 
assign N96 = ~(N48); 
assign N97 = ~(N7); 
assign N98 = ~(N27); 
assign N99 = ~(N87); 
assign N100 = ~(N8); 
assign N101 = ~(N4); 
assign N102 = ~(N88); 
assign N103 = N38 | N4; 
assign N104 = ~(N80); 
assign N105 = N53 | N6; 
assign N106 = ~(N81); 
assign N107 = ~(N84); 
assign N108 = N49 | N66; 
assign N109 = ~(N7); 
assign N110 = ~(N51); 
assign N111 = ~(N78); 
assign N112 = N18 | N76; 
assign N113 = ~(N79); 
assign N114 = ~(N16); 
assign N115 = ~(N88); 
assign N116 = ~(N17); 
assign N117 = ~(N87); 
assign N118 = N14 & N54; 
assign N119 = ~(N81); 
assign N120 = ~(N2); 
assign N121 = ~(N83); 
assign N122 = ~(N81); 
assign N123 = ~(N87); 
assign N124 = N68 & N40; 
assign N125 = ~(N41); 
assign N126 = ~(N85); 
assign N127 = ~(N53); 
assign N128 = ~(N59); 
assign N129 = N42 | N3; 
assign N130 = ~(N82); 
assign N131 = ~(N42); 
assign N132 = ~(N34); 
assign N133 = ~(N82); 
assign N134 = ~(N9); 
assign N135 = ~(N88); 
assign N136 = ~(N115); 
assign N137 = ~(N82); 
assign N138 = ~(N83); 
assign N139 = ~(N13); 
assign N140 = ~(N16); 
assign N141 = N100 & N84; 
assign N142 = N99 & N115; 
assign N143 = ~(N88); 
assign N144 = ~(N50); 
assign N145 = ~(N83); 
assign N146 = ~(N99); 
assign N147 = ~(N14); 
assign N148 = ~(N99); 
assign N149 = ~(N26); 
assign N150 = N92 | N52; 
assign N151 = ~(N84); 
assign N152 = ~(N113); 
assign N153 = ~(N127); 
assign N154 = N101 & N103; 
assign N155 = ~(N22); 
assign N156 = ~(N83); 
assign N157 = ~(N8); 
assign N158 = ~(N61); 
assign N159 = ~(N9); 
assign N160 = N74 | N122; 
assign N161 = ~(N35); 
assign N162 = ~(N89); 
assign N163 = ~(N119); 
assign N164 = ~(N78); 
assign N165 = N62 & N30; 
assign N166 = ~(N13); 
assign N167 = ~(N38); 
assign N168 = N61 | N83 | N6; 
assign N169 = ~(N86); 
assign N170 = ~(N44); 
assign N171 = ~(N56); 
assign N172 = ~(N93); 
assign N173 = ~(N102); 
assign N174 = ~(N104); 
assign N175 = ~(N121); 
assign N176 = ~(N11); 
assign N177 = ~(N16); 
assign N178 = N25 | N26 | N72; 
assign N179 = ~(N166); 
assign N180 = N19 | N51 | N151 | N159 | N174; 
assign N181 = N147 & N163; 
assign N182 = N8 | N15 | N76; 
assign N183 = N1 & N111; 
assign N184 = ~(N112); 
assign N185 = N73 & N33; 
assign N186 = N129 | N165; 
assign N187 = N27 & N81; 
assign N188 = N124 & N11; 
assign N189 = N9 & N87; 
assign N190 = N109 | N113 | N78; 
assign N191 = N148 & N169; 
assign N192 = ~(N20); 
assign N193 = N187 & N66; 
assign N194 = N7 & N71; 
assign N195 = N75 | N25; 
assign N196 = N33 | N118; 
assign N197 = N10 | N30 | N111 | N185 | N114; 
assign N198 = N161 | N30; 
assign N199 = N21 | N88; 
assign N200 = N50 & N68; 
assign N201 = N130 | N175; 
assign N202 = ~(N123); 
assign N203 = N34 & N86 & N62; 
assign N204 = ~(N89); 
assign N205 = N155 & N128; 
assign N206 = N172 | N171; 
assign N207 = N138 | N142 | N101; 
assign N208 = N6 | N131; 
assign N209 = ~(N113); 
assign N210 = ~(N141); 
assign N211 = ~(N127); 
assign N212 = ~(N7); 
assign N213 = N41 | N121 | N196 | N184; 
assign N214 = N125 | N188 | N189 | N78; 
assign N215 = N139 & N201; 
assign N216 = N52 | N66 | N182 | N165; 
assign N217 = N47 & N86; 
assign N218 = N65 | N108 | N137 | N199; 
assign N219 = ~(N196); 
assign N220 = N28 | N87 | N145 | N9; 
assign N221 = N23 & N168; 
assign N222 = N119 & N211; 
assign N223 = N135 | N160 | N170 | N162; 
assign N224 = N2 & N193 & N209; 
assign N225 = N186 | N159; 
assign N226 = N20 | N32 | N118 | N123 | N219; 
assign N227 = N149 & N198 & N219; 
assign N228 = ~(N92); 
assign N229 = N67 | N99; 
assign N230 = N59 | N95 | N143 | N144 | N191; 
assign N231 = ~(N8); 
assign N232 = ~(N212); 
assign N233 = N39 | N85 | N107 | N176 | N79; 
assign N234 = N202 & N216 & N18; 
assign N235 = N40 | N117 | N56; 
assign N236 = N16 | N88 | N133 | N107; 
assign N237 = ~(N183); 
assign N238 = ~(N222); 
assign N239 = N36 | N56 | N116 | N211; 
assign N240 = N69 & N225 & N183; 
assign N241 = N13 & N81 & N82 & N89 & N150 & N28; 
assign N242 = N4 | N233 | N53; 
assign N243 = N12 & N157 & N133; 
assign N244 = N17 | N127 | N173 | N195; 
assign N245 = N84 | N194 | N118; 
assign N246 = N90 | N206 | N218 | N220 | N231 | N36; 
assign N247 = N227 | N194; 
assign N248 = ~(N55); 
assign N249 = ~(N219); 
assign N250 = ~(N95); 
assign N251 = N94 | N175 | N199; 
assign N252 = N77 | N223; 
assign N253 = N207 & N196; 
assign N254 = ~(N54); 
assign N255 = ~(N181); 
assign N256 = N165 | N210; 
assign N257 = ~(N19); 
assign N258 = N80 & N185; 
assign N259 = N48 | N221 | N144; 
assign N260 = N131 | N178 | N142; 
assign N261 = N78 | N104 | N105 | N42; 
assign N262 = N60 & N103 & N120 & N229 & N61; 
assign N263 = N44 & N201 & N210 & N30; 
assign N264 = N190 | N203; 
assign N265 = N102 & N2; 
assign N266 = ~(N193); 
assign N267 = N251 & N186; 
assign N268 = ~(N69); 
assign N269 = ~(N147); 
assign N270 = ~(N228); 
assign N271 = N46 | N17; 
assign N272 = N255 | N202; 
assign N273 = N259 | N200; 
assign N274 = N93 & N137; 
assign N275 = ~(N214); 
assign N276 = N247 & N207; 
assign N277 = N58 & N226 & N242 & N178; 
assign N278 = N43 | N132 | N183; 
assign N279 = N249 | N176; 
assign N280 = N70 & N154; 
assign N281 = ~(N136); 
assign N282 = N228 | N218; 
assign N283 = N152 | N212 | N186; 
assign N284 = N180 | N281 | N126; 
assign N285 = N106 | N204 | N263; 
assign N286 = N91 & N171 & N268 & N84; 
assign N287 = ~(N209); 
assign N288 = N141 & N23; 
assign N289 = ~(N113); 
assign N290 = N114 & N279 & N25; 
assign N291 = N266 | N271 | N276 | N185; 
assign N292 = ~(N67); 
assign N293 = N264 & N52; 
assign N294 = N98 & N126 & N273 & N37; 
assign N295 = N122 & N169 & N197 & N256 & N261; 
assign N296 = ~(N191); 
assign N297 = N112 | N232; 
assign N298 = N153 & N183; 
assign N299 = N283 | N1; 
assign N300 = N115 & N85; 
assign N301 = ~(N2); 
assign N302 = ~(N168); 
assign N303 = ~(N163); 
assign N304 = ~(N42); 
assign N305 = ~(N205); 
assign N306 = ~(N82); 
assign N307 = ~(N232); 
assign N308 = ~(N86); 
assign N309 = ~(N144); 
assign N310 = N287 & N178; 
assign N311 = ~(N159); 
assign N312 = ~(N23); 
assign N313 = ~(N202); 
assign N314 = ~(N216); 
assign N315 = ~(N242); 
assign N316 = ~(N229); 
assign N317 = ~(N183); 
assign N318 = ~(N50); 
assign N319 = ~(N224); 
assign N320 = ~(N154); 
assign N321 = ~(N213); 
assign N322 = ~(N235); 
assign N323 = ~(N31); 
assign N324 = ~(N169); 
assign N325 = N162 & N257 & N35; 
assign N326 = N237 & N133; 
assign N327 = ~(N29); 
assign N328 = ~(N85); 
assign N329 = ~(N128); 
assign N330 = ~(N247); 
assign N331 = ~(N208); 
assign N332 = ~(N135); 
assign N333 = ~(N193); 
assign N334 = ~(N6); 
assign N335 = N110 & N196; 
assign N336 = ~(N39); 
assign N337 = ~(N195); 
assign N338 = ~(N1); 
assign N339 = ~(N184); 
assign N340 = ~(N193); 
assign N341 = ~(N211); 
assign N342 = ~(N214); 
assign N343 = N246 & N296; 
assign N344 = ~(N11); 
assign N345 = N97 | N286; 
assign N346 = ~(N96); 
assign N347 = ~(N4); 
assign N348 = N289 | N234; 
assign N349 = ~(N238); 
assign N350 = N297 & N140; 
assign N351 = ~(N193); 
assign N352 = ~(N18); 
assign N353 = ~(N262); 
assign N354 = N258 | N272; 
assign N355 = ~(N181); 
assign N356 = ~(N248); 
assign N357 = ~(N225); 
assign N358 = N195 & N41; 
assign N359 = ~(N24); 
assign N360 = ~(N78); 
assign N361 = N140 & N230; 
assign N362 = ~(N134); 
assign N363 = N267 | N216; 
assign N364 = ~(N202); 
assign N365 = ~(N139); 
assign N366 = ~(N105); 
assign N367 = ~(N91); 
assign N368 = N243 | N231; 
assign N369 = ~(N259); 
assign N370 = ~(N226); 
assign N371 = N236 | N188; 
assign N372 = ~(N89); 
assign N373 = ~(N231); 
assign N374 = ~(N223); 
assign N375 = ~(N198); 
assign N376 = ~(N65); 
assign N377 = ~(N175); 
assign N378 = ~(N186); 
assign N379 = N128 & N219 & N41; 
assign N380 = ~(N138); 
assign N381 = N277 | N180; 
assign N382 = ~(N179); 
assign N383 = ~(N338); 
assign N384 = N330 & N378 & N39; 
assign N385 = N209 | N76; 
assign N386 = N167 & N204; 
assign N387 = N333 | N218; 
assign N388 = N349 & N217; 
assign N389 = N192 & N254; 
assign N390 = ~(N252); 
assign N391 = N168 | N42; 
assign N392 = ~(N142); 
assign N393 = N278 | N300 | N61; 
assign N394 = ~(N294); 
assign N395 = N146 & N331 & N202; 
assign N396 = N260 | N302 | N340 | N165; 
assign N397 = N158 & N262 & N186; 
assign N398 = N234 | N47; 
assign N399 = N200 & N280; 
assign N400 = N274 | N228; 
assign N401 = N298 | N110; 
assign N402 = ~(N375); 
assign N403 = ~(N177); 
assign N404 = ~(N179); 
assign N405 = N164 | N66; 
assign N406 = N307 | N351 | N381 | N38; 
assign N407 = N250 | N169; 
assign N408 = N179 | N374 | N149; 
assign N409 = N373 | N121; 
assign N410 = N156 | N224; 
assign N411 = N301 & N322 & N60; 
assign N412 = ~(N199); 
assign N413 = ~(N140); 
assign N414 = N352 & N69; 
assign N415 = ~(N130); 
assign N416 = N320 | N358 | N24; 
assign N417 = N245 | N308 | N86; 
assign N418 = N345 & N208; 
assign N419 = N270 | N319 | N36; 
assign N420 = N184 & N295 & N403 & N100; 
assign N421 = ~(N48); 
assign N422 = N191 & N326 & N376 & N20; 
assign N423 = ~(N377); 
assign N424 = N230 | N288 | N327 | N338 | N188; 
assign N425 = N211 & N207; 
assign N426 = N346 & N368 & N398 & N182; 
assign N427 = N205 | N208 | N299 | N407 | N181; 
assign N428 = ~(N247); 
assign N429 = N217 & N314 & N387 & N152; 
assign N430 = ~(N272); 
assign N431 = N305 | N26; 
assign N432 = N409 | N40; 
assign N433 = ~(N222); 
assign N434 = N181 & N382 & N96; 
assign N435 = N241 & N284 & N336 & N417 & N146; 
assign N436 = N347 | N148; 
assign N437 = N290 & N356 & N366 & N115; 
assign N438 = N252 | N253 | N315 | N360 | N380 | N389 | N396 | N399; 
assign N439 = N311 & N321 & N350 & N353 & N363 & N367 & N369 & N379 & N415; 
assign N440 = N362 & N372 & N400 & N413 & N182; 
assign N441 = N213 | N304 | N306 | N316 | N365 | N408 | N414 | N423 | N437; 
assign N442 = N203 & N215 & N293 & N324 & N332 & N337 & N357 & N397 & N410; 
assign N443 = N214 | N282 | N334 | N361 | N388 | N390 | N412 | N416; 
assign N444 = ~(N25); 
assign N445 = N318 & N371 & N392 & N405; 
assign N446 = ~(N275); 
assign N447 = N335 & N344; 
assign N448 = N309 | N348; 
assign N449 = ~(N420); 
assign N450 = ~(N428); 
assign N451 = ~(N44); 
assign N452 = N419 & N434; 
assign N453 = ~(N394); 
assign N454 = ~(N430); 
assign N455 = N383 | N436; 
assign N456 = N303 | N312; 
assign N457 = N292 | N406 | N440; 
assign N458 = N385 & N433; 
assign N459 = N224 & N342 & N429 & N435; 
assign N460 = N317 | N404 | N427; 
assign N461 = N343 & N402; 
assign N462 = N244 & N325; 
assign N463 = ~(N412); 
assign N464 = ~(N235); 
assign N465 = N339 | N370 | N431 | N411; 
assign N466 = ~(N439); 
assign N467 = ~(N425); 
assign N468 = N239 | N421 | N441; 
assign N469 = ~(N392); 
assign N470 = N291 | N323 | N329; 
assign N471 = N238 & N269 & N355 & N438 & N424; 
assign N472 = N354 | N359; 
assign N473 = ~(N386); 
assign N474 = N328 & N384 & N391; 
assign N475 = N240 & N426 & N432; 
assign N476 = N265 | N395 | N443; 
assign N477 = N313 & N364 & N401 & N418; 
assign N478 = ~(N393); 
assign N479 = N341 & N422 & N439 & N442; 
assign N480 = ~(N285); 
assign N481 = ~(N310); 
endmodule
