module Depth_10_20_Nodes_200_400_S009 (N1, N2, N3, N4, N5, N6, N7, N8, N275, N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286, N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297, N298, N299, N300);

input N1; 
input N2; 
input N3; 
input N4; 
input N5; 
input N6; 
input N7; 
input N8; 

output N275; 
output N276; 
output N277; 
output N278; 
output N279; 
output N280; 
output N281; 
output N282; 
output N283; 
output N284; 
output N285; 
output N286; 
output N287; 
output N288; 
output N289; 
output N290; 
output N291; 
output N292; 
output N293; 
output N294; 
output N295; 
output N296; 
output N297; 
output N298; 
output N299; 
output N300; 

wire N9; 
wire N10; 
wire N11; 
wire N12; 
wire N13; 
wire N14; 
wire N15; 
wire N16; 
wire N17; 
wire N18; 
wire N19; 
wire N20; 
wire N21; 
wire N22; 
wire N23; 
wire N24; 
wire N25; 
wire N26; 
wire N27; 
wire N28; 
wire N29; 
wire N30; 
wire N31; 
wire N32; 
wire N33; 
wire N34; 
wire N35; 
wire N36; 
wire N37; 
wire N38; 
wire N39; 
wire N40; 
wire N41; 
wire N42; 
wire N43; 
wire N44; 
wire N45; 
wire N46; 
wire N47; 
wire N48; 
wire N49; 
wire N50; 
wire N51; 
wire N52; 
wire N53; 
wire N54; 
wire N55; 
wire N56; 
wire N57; 
wire N58; 
wire N59; 
wire N60; 
wire N61; 
wire N62; 
wire N63; 
wire N64; 
wire N65; 
wire N66; 
wire N67; 
wire N68; 
wire N69; 
wire N70; 
wire N71; 
wire N72; 
wire N73; 
wire N74; 
wire N75; 
wire N76; 
wire N77; 
wire N78; 
wire N79; 
wire N80; 
wire N81; 
wire N82; 
wire N83; 
wire N84; 
wire N85; 
wire N86; 
wire N87; 
wire N88; 
wire N89; 
wire N90; 
wire N91; 
wire N92; 
wire N93; 
wire N94; 
wire N95; 
wire N96; 
wire N97; 
wire N98; 
wire N99; 
wire N100; 
wire N101; 
wire N102; 
wire N103; 
wire N104; 
wire N105; 
wire N106; 
wire N107; 
wire N108; 
wire N109; 
wire N110; 
wire N111; 
wire N112; 
wire N113; 
wire N114; 
wire N115; 
wire N116; 
wire N117; 
wire N118; 
wire N119; 
wire N120; 
wire N121; 
wire N122; 
wire N123; 
wire N124; 
wire N125; 
wire N126; 
wire N127; 
wire N128; 
wire N129; 
wire N130; 
wire N131; 
wire N132; 
wire N133; 
wire N134; 
wire N135; 
wire N136; 
wire N137; 
wire N138; 
wire N139; 
wire N140; 
wire N141; 
wire N142; 
wire N143; 
wire N144; 
wire N145; 
wire N146; 
wire N147; 
wire N148; 
wire N149; 
wire N150; 
wire N151; 
wire N152; 
wire N153; 
wire N154; 
wire N155; 
wire N156; 
wire N157; 
wire N158; 
wire N159; 
wire N160; 
wire N161; 
wire N162; 
wire N163; 
wire N164; 
wire N165; 
wire N166; 
wire N167; 
wire N168; 
wire N169; 
wire N170; 
wire N171; 
wire N172; 
wire N173; 
wire N174; 
wire N175; 
wire N176; 
wire N177; 
wire N178; 
wire N179; 
wire N180; 
wire N181; 
wire N182; 
wire N183; 
wire N184; 
wire N185; 
wire N186; 
wire N187; 
wire N188; 
wire N189; 
wire N190; 
wire N191; 
wire N192; 
wire N193; 
wire N194; 
wire N195; 
wire N196; 
wire N197; 
wire N198; 
wire N199; 
wire N200; 
wire N201; 
wire N202; 
wire N203; 
wire N204; 
wire N205; 
wire N206; 
wire N207; 
wire N208; 
wire N209; 
wire N210; 
wire N211; 
wire N212; 
wire N213; 
wire N214; 
wire N215; 
wire N216; 
wire N217; 
wire N218; 
wire N219; 
wire N220; 
wire N221; 
wire N222; 
wire N223; 
wire N224; 
wire N225; 
wire N226; 
wire N227; 
wire N228; 
wire N229; 
wire N230; 
wire N231; 
wire N232; 
wire N233; 
wire N234; 
wire N235; 
wire N236; 
wire N237; 
wire N238; 
wire N239; 
wire N240; 
wire N241; 
wire N242; 
wire N243; 
wire N244; 
wire N245; 
wire N246; 
wire N247; 
wire N248; 
wire N249; 
wire N250; 
wire N251; 
wire N252; 
wire N253; 
wire N254; 
wire N255; 
wire N256; 
wire N257; 
wire N258; 
wire N259; 
wire N260; 
wire N261; 
wire N262; 
wire N263; 
wire N264; 
wire N265; 
wire N266; 
wire N267; 
wire N268; 
wire N269; 
wire N270; 
wire N271; 
wire N272; 
wire N273; 
wire N274; 

assign N9 = ~(N4); 
assign N10 = ~(N4); 
assign N11 = ~(N5); 
assign N12 = ~(N8); 
assign N13 = ~(N3); 
assign N14 = ~(N2); 
assign N15 = ~(N6); 
assign N16 = ~(N1); 
assign N17 = ~(N8); 
assign N18 = ~(N7); 
assign N19 = ~(N5); 
assign N20 = ~(N8); 
assign N21 = ~(N4); 
assign N22 = ~(N3); 
assign N23 = ~(N5); 
assign N24 = ~(N2); 
assign N25 = ~(N2); 
assign N26 = ~(N7); 
assign N27 = ~(N6); 
assign N28 = ~(N27); 
assign N29 = ~(N20); 
assign N30 = N1 | N5; 
assign N31 = ~(N2); 
assign N32 = ~(N26); 
assign N33 = ~(N22); 
assign N34 = ~(N19); 
assign N35 = N18 & N23; 
assign N36 = ~(N6); 
assign N37 = ~(N6); 
assign N38 = ~(N13); 
assign N39 = ~(N28); 
assign N40 = ~(N37); 
assign N41 = ~(N21); 
assign N42 = ~(N28); 
assign N43 = ~(N32); 
assign N44 = ~(N8); 
assign N45 = ~(N13); 
assign N46 = ~(N29); 
assign N47 = ~(N34); 
assign N48 = ~(N38); 
assign N49 = N38 | N9; 
assign N50 = ~(N12); 
assign N51 = N32 | N10; 
assign N52 = ~(N26); 
assign N53 = N10 | N29 | N15; 
assign N54 = ~(N7); 
assign N55 = ~(N28); 
assign N56 = ~(N42); 
assign N57 = ~(N51); 
assign N58 = ~(N36); 
assign N59 = ~(N40); 
assign N60 = ~(N44); 
assign N61 = ~(N12); 
assign N62 = N19 | N3; 
assign N63 = ~(N51); 
assign N64 = ~(N19); 
assign N65 = ~(N30); 
assign N66 = ~(N40); 
assign N67 = ~(N22); 
assign N68 = ~(N39); 
assign N69 = ~(N50); 
assign N70 = ~(N14); 
assign N71 = ~(N24); 
assign N72 = ~(N7); 
assign N73 = ~(N35); 
assign N74 = ~(N27); 
assign N75 = ~(N7); 
assign N76 = ~(N16); 
assign N77 = ~(N33); 
assign N78 = ~(N52); 
assign N79 = ~(N36); 
assign N80 = ~(N15); 
assign N81 = ~(N17); 
assign N82 = ~(N38); 
assign N83 = N6 | N47; 
assign N84 = ~(N5); 
assign N85 = ~(N42); 
assign N86 = ~(N53); 
assign N87 = ~(N45); 
assign N88 = ~(N48); 
assign N89 = ~(N51); 
assign N90 = ~(N6); 
assign N91 = ~(N28); 
assign N92 = ~(N15); 
assign N93 = ~(N11); 
assign N94 = ~(N36); 
assign N95 = ~(N13); 
assign N96 = ~(N22); 
assign N97 = ~(N42); 
assign N98 = ~(N32); 
assign N99 = ~(N26); 
assign N100 = ~(N24); 
assign N101 = ~(N33); 
assign N102 = ~(N34); 
assign N103 = ~(N44); 
assign N104 = ~(N18); 
assign N105 = ~(N33); 
assign N106 = ~(N4); 
assign N107 = ~(N41); 
assign N108 = ~(N24); 
assign N109 = ~(N39); 
assign N110 = N2 & N33 & N45; 
assign N111 = ~(N34); 
assign N112 = ~(N40); 
assign N113 = ~(N47); 
assign N114 = ~(N20); 
assign N115 = ~(N52); 
assign N116 = ~(N20); 
assign N117 = ~(N45); 
assign N118 = ~(N31); 
assign N119 = ~(N36); 
assign N120 = N69 & N32; 
assign N121 = ~(N27); 
assign N122 = ~(N42); 
assign N123 = ~(N22); 
assign N124 = N57 | N19; 
assign N125 = ~(N86); 
assign N126 = ~(N28); 
assign N127 = ~(N114); 
assign N128 = N3 & N95; 
assign N129 = ~(N51); 
assign N130 = ~(N48); 
assign N131 = ~(N34); 
assign N132 = N76 & N31; 
assign N133 = N56 & N94 & N108; 
assign N134 = ~(N79); 
assign N135 = ~(N3); 
assign N136 = ~(N16); 
assign N137 = N41 | N29; 
assign N138 = N97 & N50; 
assign N139 = N78 & N19; 
assign N140 = N17 & N80 & N37; 
assign N141 = N9 | N39; 
assign N142 = ~(N35); 
assign N143 = N63 | N46; 
assign N144 = N42 | N53 | N13; 
assign N145 = N102 | N31; 
assign N146 = ~(N137); 
assign N147 = ~(N123); 
assign N148 = N36 & N45 & N129; 
assign N149 = N4 & N27 & N68 & N113; 
assign N150 = ~(N114); 
assign N151 = ~(N41); 
assign N152 = ~(N126); 
assign N153 = N14 | N101 | N107 | N131 | N50; 
assign N154 = N140 | N13; 
assign N155 = N21 | N58 | N43; 
assign N156 = N51 | N118 | N126 | N136; 
assign N157 = N133 & N121; 
assign N158 = ~(N15); 
assign N159 = N117 | N1; 
assign N160 = ~(N33); 
assign N161 = ~(N34); 
assign N162 = N66 | N154; 
assign N163 = ~(N72); 
assign N164 = ~(N1); 
assign N165 = ~(N30); 
assign N166 = ~(N153); 
assign N167 = N39 & N144; 
assign N168 = N104 | N49; 
assign N169 = N28 | N158; 
assign N170 = ~(N93); 
assign N171 = N37 & N59 & N91; 
assign N172 = ~(N7); 
assign N173 = ~(N52); 
assign N174 = N87 | N108 | N45; 
assign N175 = N99 & N139 & N147 & N122; 
assign N176 = N22 | N132 | N50; 
assign N177 = N116 & N107; 
assign N178 = ~(N21); 
assign N179 = N125 & N130 & N144; 
assign N180 = ~(N32); 
assign N181 = N24 | N100 | N106 | N143 | N118; 
assign N182 = N153 | N171 | N180; 
assign N183 = N20 | N65 | N34; 
assign N184 = N11 | N23 | N31 | N89 | N158 | N176; 
assign N185 = N8 | N35 | N48 | N64 | N84 | N88 | N152 | N165; 
assign N186 = N163 & N18; 
assign N187 = ~(N153); 
assign N188 = N142 | N27; 
assign N189 = N81 & N154 & N20; 
assign N190 = N67 | N86 | N98 | N128 | N141 | N160 | N99; 
assign N191 = ~(N160); 
assign N192 = N151 & N174 & N35; 
assign N193 = N122 & N152; 
assign N194 = N5 & N12 & N129 & N163; 
assign N195 = N43 & N138 & N148 & N174; 
assign N196 = N16 | N49; 
assign N197 = N74 & N161 & N178 & N189 & N122; 
assign N198 = ~(N161); 
assign N199 = ~(N152); 
assign N200 = ~(N64); 
assign N201 = N47 | N50 | N135 | N85; 
assign N202 = ~(N157); 
assign N203 = ~(N110); 
assign N204 = ~(N181); 
assign N205 = N155 & N168 & N185 & N182; 
assign N206 = N188 & N30; 
assign N207 = ~(N115); 
assign N208 = N167 & N144; 
assign N209 = N40 & N166 & N177; 
assign N210 = N13 | N134 | N52; 
assign N211 = N25 | N26; 
assign N212 = N46 | N90; 
assign N213 = N79 | N82 | N83 | N111 | N127 | N164 | N190 | N84; 
assign N214 = N44 | N72 | N194 | N70; 
assign N215 = N30 & N55 & N60 & N62 & N105 & N109 & N181 & N182; 
assign N216 = N54 | N61 | N93 | N187 | N191 | N204 | N181; 
assign N217 = ~(N44); 
assign N218 = ~(N112); 
assign N219 = N73 & N119 & N149 & N200 & N207; 
assign N220 = N70 | N115 | N121 | N41; 
assign N221 = N183 & N211 & N118; 
assign N222 = N173 | N177 | N196; 
assign N223 = N71 & N146; 
assign N224 = ~(N184); 
assign N225 = ~(N182); 
assign N226 = ~(N91); 
assign N227 = N103 & N132; 
assign N228 = N75 | N203 | N166; 
assign N229 = N92 & N157 & N170 & N209 & N137; 
assign N230 = ~(N176); 
assign N231 = N208 | N39; 
assign N232 = ~(N53); 
assign N233 = N85 | N14; 
assign N234 = N206 & N183; 
assign N235 = N175 & N186 & N112; 
assign N236 = N150 & N93; 
assign N237 = ~(N145); 
assign N238 = ~(N32); 
assign N239 = ~(N51); 
assign N240 = N77 | N216 | N124; 
assign N241 = N212 | N54; 
assign N242 = N96 | N156 | N214 | N172; 
assign N243 = N124 & N165 & N185; 
assign N244 = N241 & N31; 
assign N245 = N197 | N199 | N219 | N130; 
assign N246 = ~(N145); 
assign N247 = N198 & N202 & N230 & N239 & N242 & N125; 
assign N248 = ~(N109); 
assign N249 = ~(N148); 
assign N250 = N233 | N179; 
assign N251 = N146 & N210 & N238 & N176; 
assign N252 = ~(N40); 
assign N253 = N136 | N10; 
assign N254 = N120 & N227 & N14; 
assign N255 = N159 | N180 | N193 | N222; 
assign N256 = N249 & N176; 
assign N257 = N250 | N129; 
assign N258 = ~(N185); 
assign N259 = N220 & N164; 
assign N260 = ~(N31); 
assign N261 = N232 | N155; 
assign N262 = ~(N235); 
assign N263 = N228 | N248 | N130; 
assign N264 = ~(N149); 
assign N265 = ~(N154); 
assign N266 = ~(N244); 
assign N267 = N195 & N46; 
assign N268 = N221 & N125; 
assign N269 = N179 & N237; 
assign N270 = ~(N168); 
assign N271 = N252 | N183; 
assign N272 = N229 & N182; 
assign N273 = N225 & N148; 
assign N274 = ~(N169); 
assign N275 = N240 | N243 | N266; 
assign N276 = ~(N231); 
assign N277 = ~(N274); 
assign N278 = ~(N46); 
assign N279 = ~(N236); 
assign N280 = N205 | N258; 
assign N281 = N215 & N251 & N273; 
assign N282 = N162 | N245; 
assign N283 = ~(N224); 
assign N284 = ~(N260); 
assign N285 = N253 & N259; 
assign N286 = ~(N268); 
assign N287 = ~(N261); 
assign N288 = ~(N247); 
assign N289 = ~(N99); 
assign N290 = N192 | N255 | N257; 
assign N291 = N223 & N256 & N264; 
assign N292 = N218 & N226 & N269; 
assign N293 = N184 & N267 & N270 & N272; 
assign N294 = ~(N260); 
assign N295 = ~(N265); 
assign N296 = N201 | N234 | N262; 
assign N297 = N213 & N254; 
assign N298 = ~(N172); 
assign N299 = ~(N263); 
assign N300 = N217 & N246 & N265 & N271; 
endmodule
