module Depth_10_20_Nodes_200_400_S008 (N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N356, N357, N358, N359, N360, N361, N362, N363, N364, N365, N366, N367, N368, N369, N370, N371, N372, N373, N374, N375, N376, N377, N378);

input N1; 
input N2; 
input N3; 
input N4; 
input N5; 
input N6; 
input N7; 
input N8; 
input N9; 
input N10; 
input N11; 
input N12; 
input N13; 

output N356; 
output N357; 
output N358; 
output N359; 
output N360; 
output N361; 
output N362; 
output N363; 
output N364; 
output N365; 
output N366; 
output N367; 
output N368; 
output N369; 
output N370; 
output N371; 
output N372; 
output N373; 
output N374; 
output N375; 
output N376; 
output N377; 
output N378; 

wire N14; 
wire N15; 
wire N16; 
wire N17; 
wire N18; 
wire N19; 
wire N20; 
wire N21; 
wire N22; 
wire N23; 
wire N24; 
wire N25; 
wire N26; 
wire N27; 
wire N28; 
wire N29; 
wire N30; 
wire N31; 
wire N32; 
wire N33; 
wire N34; 
wire N35; 
wire N36; 
wire N37; 
wire N38; 
wire N39; 
wire N40; 
wire N41; 
wire N42; 
wire N43; 
wire N44; 
wire N45; 
wire N46; 
wire N47; 
wire N48; 
wire N49; 
wire N50; 
wire N51; 
wire N52; 
wire N53; 
wire N54; 
wire N55; 
wire N56; 
wire N57; 
wire N58; 
wire N59; 
wire N60; 
wire N61; 
wire N62; 
wire N63; 
wire N64; 
wire N65; 
wire N66; 
wire N67; 
wire N68; 
wire N69; 
wire N70; 
wire N71; 
wire N72; 
wire N73; 
wire N74; 
wire N75; 
wire N76; 
wire N77; 
wire N78; 
wire N79; 
wire N80; 
wire N81; 
wire N82; 
wire N83; 
wire N84; 
wire N85; 
wire N86; 
wire N87; 
wire N88; 
wire N89; 
wire N90; 
wire N91; 
wire N92; 
wire N93; 
wire N94; 
wire N95; 
wire N96; 
wire N97; 
wire N98; 
wire N99; 
wire N100; 
wire N101; 
wire N102; 
wire N103; 
wire N104; 
wire N105; 
wire N106; 
wire N107; 
wire N108; 
wire N109; 
wire N110; 
wire N111; 
wire N112; 
wire N113; 
wire N114; 
wire N115; 
wire N116; 
wire N117; 
wire N118; 
wire N119; 
wire N120; 
wire N121; 
wire N122; 
wire N123; 
wire N124; 
wire N125; 
wire N126; 
wire N127; 
wire N128; 
wire N129; 
wire N130; 
wire N131; 
wire N132; 
wire N133; 
wire N134; 
wire N135; 
wire N136; 
wire N137; 
wire N138; 
wire N139; 
wire N140; 
wire N141; 
wire N142; 
wire N143; 
wire N144; 
wire N145; 
wire N146; 
wire N147; 
wire N148; 
wire N149; 
wire N150; 
wire N151; 
wire N152; 
wire N153; 
wire N154; 
wire N155; 
wire N156; 
wire N157; 
wire N158; 
wire N159; 
wire N160; 
wire N161; 
wire N162; 
wire N163; 
wire N164; 
wire N165; 
wire N166; 
wire N167; 
wire N168; 
wire N169; 
wire N170; 
wire N171; 
wire N172; 
wire N173; 
wire N174; 
wire N175; 
wire N176; 
wire N177; 
wire N178; 
wire N179; 
wire N180; 
wire N181; 
wire N182; 
wire N183; 
wire N184; 
wire N185; 
wire N186; 
wire N187; 
wire N188; 
wire N189; 
wire N190; 
wire N191; 
wire N192; 
wire N193; 
wire N194; 
wire N195; 
wire N196; 
wire N197; 
wire N198; 
wire N199; 
wire N200; 
wire N201; 
wire N202; 
wire N203; 
wire N204; 
wire N205; 
wire N206; 
wire N207; 
wire N208; 
wire N209; 
wire N210; 
wire N211; 
wire N212; 
wire N213; 
wire N214; 
wire N215; 
wire N216; 
wire N217; 
wire N218; 
wire N219; 
wire N220; 
wire N221; 
wire N222; 
wire N223; 
wire N224; 
wire N225; 
wire N226; 
wire N227; 
wire N228; 
wire N229; 
wire N230; 
wire N231; 
wire N232; 
wire N233; 
wire N234; 
wire N235; 
wire N236; 
wire N237; 
wire N238; 
wire N239; 
wire N240; 
wire N241; 
wire N242; 
wire N243; 
wire N244; 
wire N245; 
wire N246; 
wire N247; 
wire N248; 
wire N249; 
wire N250; 
wire N251; 
wire N252; 
wire N253; 
wire N254; 
wire N255; 
wire N256; 
wire N257; 
wire N258; 
wire N259; 
wire N260; 
wire N261; 
wire N262; 
wire N263; 
wire N264; 
wire N265; 
wire N266; 
wire N267; 
wire N268; 
wire N269; 
wire N270; 
wire N271; 
wire N272; 
wire N273; 
wire N274; 
wire N275; 
wire N276; 
wire N277; 
wire N278; 
wire N279; 
wire N280; 
wire N281; 
wire N282; 
wire N283; 
wire N284; 
wire N285; 
wire N286; 
wire N287; 
wire N288; 
wire N289; 
wire N290; 
wire N291; 
wire N292; 
wire N293; 
wire N294; 
wire N295; 
wire N296; 
wire N297; 
wire N298; 
wire N299; 
wire N300; 
wire N301; 
wire N302; 
wire N303; 
wire N304; 
wire N305; 
wire N306; 
wire N307; 
wire N308; 
wire N309; 
wire N310; 
wire N311; 
wire N312; 
wire N313; 
wire N314; 
wire N315; 
wire N316; 
wire N317; 
wire N318; 
wire N319; 
wire N320; 
wire N321; 
wire N322; 
wire N323; 
wire N324; 
wire N325; 
wire N326; 
wire N327; 
wire N328; 
wire N329; 
wire N330; 
wire N331; 
wire N332; 
wire N333; 
wire N334; 
wire N335; 
wire N336; 
wire N337; 
wire N338; 
wire N339; 
wire N340; 
wire N341; 
wire N342; 
wire N343; 
wire N344; 
wire N345; 
wire N346; 
wire N347; 
wire N348; 
wire N349; 
wire N350; 
wire N351; 
wire N352; 
wire N353; 
wire N354; 
wire N355; 

assign N14 = ~(N2); 
assign N15 = ~(N6); 
assign N16 = ~(N6); 
assign N17 = ~(N6); 
assign N18 = ~(N11); 
assign N19 = ~(N11); 
assign N20 = ~(N5); 
assign N21 = ~(N10); 
assign N22 = ~(N2); 
assign N23 = ~(N9); 
assign N24 = ~(N6); 
assign N25 = ~(N7); 
assign N26 = ~(N9); 
assign N27 = ~(N4); 
assign N28 = ~(N1); 
assign N29 = ~(N1); 
assign N30 = ~(N1); 
assign N31 = ~(N13); 
assign N32 = N5 | N10; 
assign N33 = ~(N4); 
assign N34 = ~(N3); 
assign N35 = ~(N1); 
assign N36 = ~(N8); 
assign N37 = ~(N3); 
assign N38 = ~(N12); 
assign N39 = ~(N10); 
assign N40 = ~(N12); 
assign N41 = ~(N13); 
assign N42 = ~(N4); 
assign N43 = ~(N3); 
assign N44 = ~(N2); 
assign N45 = ~(N3); 
assign N46 = ~(N7); 
assign N47 = ~(N34); 
assign N48 = ~(N13); 
assign N49 = ~(N25); 
assign N50 = ~(N42); 
assign N51 = ~(N40); 
assign N52 = ~(N31); 
assign N53 = ~(N4); 
assign N54 = N31 & N13; 
assign N55 = ~(N18); 
assign N56 = ~(N31); 
assign N57 = ~(N23); 
assign N58 = ~(N23); 
assign N59 = N25 & N4; 
assign N60 = ~(N39); 
assign N61 = ~(N8); 
assign N62 = ~(N46); 
assign N63 = ~(N8); 
assign N64 = N13 | N8; 
assign N65 = ~(N11); 
assign N66 = N10 & N17; 
assign N67 = N34 & N28; 
assign N68 = ~(N8); 
assign N69 = N28 & N35; 
assign N70 = ~(N10); 
assign N71 = ~(N45); 
assign N72 = ~(N16); 
assign N73 = ~(N36); 
assign N74 = ~(N5); 
assign N75 = ~(N33); 
assign N76 = ~(N23); 
assign N77 = ~(N30); 
assign N78 = ~(N16); 
assign N79 = ~(N46); 
assign N80 = ~(N9); 
assign N81 = ~(N5); 
assign N82 = ~(N17); 
assign N83 = N40 & N53 & N71; 
assign N84 = N55 & N77; 
assign N85 = N7 | N12; 
assign N86 = N62 & N60; 
assign N87 = ~(N75); 
assign N88 = N75 | N70; 
assign N89 = N61 | N22; 
assign N90 = N65 & N23; 
assign N91 = ~(N18); 
assign N92 = N11 & N19 & N5; 
assign N93 = ~(N66); 
assign N94 = N84 | N89; 
assign N95 = ~(N88); 
assign N96 = ~(N43); 
assign N97 = N27 | N79 | N41; 
assign N98 = ~(N20); 
assign N99 = ~(N90); 
assign N100 = N70 | N75; 
assign N101 = ~(N54); 
assign N102 = N24 | N35; 
assign N103 = ~(N87); 
assign N104 = N16 & N62; 
assign N105 = ~(N50); 
assign N106 = ~(N88); 
assign N107 = N22 | N9; 
assign N108 = ~(N22); 
assign N109 = N33 | N42 | N26; 
assign N110 = ~(N39); 
assign N111 = ~(N82); 
assign N112 = ~(N56); 
assign N113 = N2 & N39 & N86; 
assign N114 = ~(N35); 
assign N115 = ~(N59); 
assign N116 = ~(N74); 
assign N117 = N46 & N92; 
assign N118 = ~(N91); 
assign N119 = ~(N12); 
assign N120 = ~(N63); 
assign N121 = N81 | N42; 
assign N122 = ~(N12); 
assign N123 = N86 | N17; 
assign N124 = ~(N74); 
assign N125 = N43 | N28; 
assign N126 = ~(N34); 
assign N127 = N45 | N88; 
assign N128 = N32 & N48 & N71; 
assign N129 = ~(N70); 
assign N130 = N3 & N92; 
assign N131 = ~(N56); 
assign N132 = N4 & N68 & N115 & N63; 
assign N133 = ~(N121); 
assign N134 = ~(N30); 
assign N135 = ~(N111); 
assign N136 = ~(N120); 
assign N137 = N49 & N95; 
assign N138 = ~(N88); 
assign N139 = ~(N7); 
assign N140 = ~(N81); 
assign N141 = ~(N15); 
assign N142 = N63 & N72; 
assign N143 = N64 & N35; 
assign N144 = ~(N21); 
assign N145 = N9 & N108 & N103; 
assign N146 = ~(N70); 
assign N147 = ~(N84); 
assign N148 = N57 & N119; 
assign N149 = ~(N2); 
assign N150 = N103 & N44; 
assign N151 = N122 & N39; 
assign N152 = N1 | N106 | N65; 
assign N153 = ~(N59); 
assign N154 = N6 & N90 & N112; 
assign N155 = ~(N114); 
assign N156 = N76 | N83; 
assign N157 = ~(N72); 
assign N158 = ~(N42); 
assign N159 = N12 | N91; 
assign N160 = ~(N110); 
assign N161 = ~(N82); 
assign N162 = N20 & N37; 
assign N163 = ~(N97); 
assign N164 = ~(N83); 
assign N165 = N113 & N82; 
assign N166 = N14 | N89; 
assign N167 = ~(N37); 
assign N168 = N21 & N92; 
assign N169 = N29 & N131 & N142; 
assign N170 = N44 & N80 & N89 & N127 & N129; 
assign N171 = N26 & N126 & N141; 
assign N172 = N59 | N95 | N47; 
assign N173 = ~(N166); 
assign N174 = N74 | N71; 
assign N175 = ~(N64); 
assign N176 = N60 | N78 | N89; 
assign N177 = N134 & N113; 
assign N178 = ~(N105); 
assign N179 = N116 & N92; 
assign N180 = N124 | N137 | N147 | N168; 
assign N181 = N135 | N42; 
assign N182 = N82 & N151 & N67; 
assign N183 = N105 | N136 | N27; 
assign N184 = N125 & N93; 
assign N185 = N23 | N86; 
assign N186 = N66 | N94 | N102 | N51; 
assign N187 = ~(N44); 
assign N188 = ~(N44); 
assign N189 = ~(N142); 
assign N190 = ~(N83); 
assign N191 = N87 | N142; 
assign N192 = N88 | N100; 
assign N193 = ~(N2); 
assign N194 = N15 & N83; 
assign N195 = N93 | N51; 
assign N196 = N18 & N11; 
assign N197 = N56 | N158 | N31; 
assign N198 = N38 & N140; 
assign N199 = N143 & N165 & N173 & N33; 
assign N200 = N99 & N130 & N132 & N170 & N89; 
assign N201 = N107 & N38; 
assign N202 = ~(N141); 
assign N203 = N41 & N160; 
assign N204 = ~(N164); 
assign N205 = ~(N82); 
assign N206 = ~(N115); 
assign N207 = ~(N167); 
assign N208 = N35 | N139 | N101; 
assign N209 = ~(N15); 
assign N210 = N146 | N91; 
assign N211 = ~(N148); 
assign N212 = ~(N154); 
assign N213 = ~(N162); 
assign N214 = N97 | N100; 
assign N215 = N100 | N175; 
assign N216 = N67 | N111 | N135; 
assign N217 = N191 | N26; 
assign N218 = N51 | N72 | N58; 
assign N219 = ~(N17); 
assign N220 = ~(N113); 
assign N221 = N58 & N125; 
assign N222 = N52 | N154; 
assign N223 = ~(N166); 
assign N224 = N69 & N118 & N179 & N86; 
assign N225 = ~(N87); 
assign N226 = ~(N64); 
assign N227 = ~(N24); 
assign N228 = N71 & N54; 
assign N229 = N140 & N195 & N116; 
assign N230 = ~(N132); 
assign N231 = N206 & N132; 
assign N232 = N54 & N152; 
assign N233 = ~(N199); 
assign N234 = N73 | N117 | N214 | N63; 
assign N235 = ~(N165); 
assign N236 = N186 & N128; 
assign N237 = ~(N119); 
assign N238 = N92 & N85; 
assign N239 = ~(N163); 
assign N240 = ~(N90); 
assign N241 = N47 | N103; 
assign N242 = N193 & N58; 
assign N243 = ~(N163); 
assign N244 = N101 | N180 | N113; 
assign N245 = N169 & N188 & N219; 
assign N246 = N128 & N197 & N218; 
assign N247 = N112 | N121 | N236 | N87; 
assign N248 = N119 & N167 & N106; 
assign N249 = N133 & N145 & N19; 
assign N250 = N98 | N123 | N229 | N165; 
assign N251 = N150 | N166 | N204; 
assign N252 = N185 | N139; 
assign N253 = ~(N121); 
assign N254 = N159 | N174 | N130; 
assign N255 = N203 | N20; 
assign N256 = ~(N59); 
assign N257 = ~(N163); 
assign N258 = ~(N167); 
assign N259 = N162 & N7; 
assign N260 = N104 | N114 | N152 | N123; 
assign N261 = ~(N60); 
assign N262 = ~(N63); 
assign N263 = N222 | N164; 
assign N264 = N171 | N225 | N107; 
assign N265 = N85 | N149 | N167; 
assign N266 = N148 | N189 | N232 | N39; 
assign N267 = ~(N76); 
assign N268 = N178 | N200 | N163; 
assign N269 = N156 & N192 & N241 & N93; 
assign N270 = N217 & N258 & N113; 
assign N271 = N240 | N127; 
assign N272 = ~(N35); 
assign N273 = N211 | N251 | N37; 
assign N274 = N96 | N164 | N239 | N249 | N91; 
assign N275 = N155 & N82; 
assign N276 = ~(N144); 
assign N277 = N110 | N181 | N233 | N244 | N117; 
assign N278 = N160 & N69; 
assign N279 = N109 & N129 & N27; 
assign N280 = N153 & N254 & N66; 
assign N281 = ~(N168); 
assign N282 = ~(N140); 
assign N283 = ~(N25); 
assign N284 = N207 | N36; 
assign N285 = N157 | N124; 
assign N286 = ~(N219); 
assign N287 = ~(N182); 
assign N288 = ~(N44); 
assign N289 = N262 | N90; 
assign N290 = N212 | N126; 
assign N291 = ~(N87); 
assign N292 = ~(N39); 
assign N293 = N227 | N272; 
assign N294 = N279 & N98; 
assign N295 = N242 | N59; 
assign N296 = ~(N31); 
assign N297 = N199 | N257 | N162; 
assign N298 = ~(N158); 
assign N299 = N215 | N24; 
assign N300 = ~(N129); 
assign N301 = ~(N156); 
assign N302 = ~(N173); 
assign N303 = N228 | N265; 
assign N304 = ~(N161); 
assign N305 = ~(N79); 
assign N306 = ~(N230); 
assign N307 = ~(N95); 
assign N308 = N275 | N94; 
assign N309 = N201 | N33; 
assign N310 = ~(N117); 
assign N311 = ~(N221); 
assign N312 = N246 & N131; 
assign N313 = ~(N15); 
assign N314 = ~(N126); 
assign N315 = N138 | N176 | N94; 
assign N316 = ~(N68); 
assign N317 = N220 & N136; 
assign N318 = ~(N57); 
assign N319 = ~(N84); 
assign N320 = N177 & N105; 
assign N321 = ~(N169); 
assign N322 = ~(N30); 
assign N323 = N290 | N67; 
assign N324 = ~(N213); 
assign N325 = N198 & N284 & N305; 
assign N326 = N184 | N264 | N110; 
assign N327 = N263 & N273 & N73; 
assign N328 = N190 & N234 & N289; 
assign N329 = N224 | N247 | N274; 
assign N330 = N243 & N319 & N141; 
assign N331 = ~(N48); 
assign N332 = N276 | N298 | N51; 
assign N333 = N287 & N29; 
assign N334 = N237 & N261 & N90; 
assign N335 = N194 | N252 | N288 | N293 | N108; 
assign N336 = N256 | N301 | N118; 
assign N337 = N172 & N226 & N300 & N311 & N159; 
assign N338 = N208 & N285; 
assign N339 = N216 & N231 & N122; 
assign N340 = N196 & N209; 
assign N341 = N202 | N210 | N296 | N316; 
assign N342 = ~(N103); 
assign N343 = N283 | N328 | N330; 
assign N344 = ~(N277); 
assign N345 = N187 & N248 & N286 & N302; 
assign N346 = ~(N266); 
assign N347 = N259 | N280 | N318 | N338; 
assign N348 = N307 & N84; 
assign N349 = N291 & N303 & N313 & N329 & N155; 
assign N350 = N183 & N235 & N268 & N295 & N332 & N122; 
assign N351 = N223 & N34; 
assign N352 = N255 | N118; 
assign N353 = N309 & N166; 
assign N354 = N294 & N323; 
assign N355 = N205 | N250 | N158; 
assign N356 = N312 | N315 | N343 | N350 | N355; 
assign N357 = N253 | N325 | N348; 
assign N358 = N270 | N345 | N353; 
assign N359 = N266 & N322 & N340; 
assign N360 = N281 | N306 | N334 | N336 | N339; 
assign N361 = N326 | N333 | N346; 
assign N362 = N297 & N314; 
assign N363 = N269 | N282 | N347; 
assign N364 = ~(N297); 
assign N365 = ~(N28); 
assign N366 = ~(N331); 
assign N367 = N292 | N321 | N351; 
assign N368 = N317 | N341; 
assign N369 = N260 | N342; 
assign N370 = N278 & N299; 
assign N371 = N267 | N310 | N354; 
assign N372 = ~(N92); 
assign N373 = N245 & N304 & N335; 
assign N374 = N238 | N324; 
assign N375 = N308 | N337; 
assign N376 = ~(N320); 
assign N377 = N327 & N349; 
assign N378 = N271 | N344 | N352; 
endmodule
