module Depth_10_20_Nodes_200_400_S000 (N1, N2, N3, N4, N5, N6, N415, N416, N417, N418, N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429, N430, N431, N432, N433, N434, N435, N436, N437, N438, N439, N440, N441, N442, N443, N444, N445, N446, N447, N448, N449, N450, N451, N452, N453, N454, N455, N456, N457, N458, N459, N460, N461, N462, N463, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473, N474, N475, N476, N477);

input N1; 
input N2; 
input N3; 
input N4; 
input N5; 
input N6; 

output N415; 
output N416; 
output N417; 
output N418; 
output N419; 
output N420; 
output N421; 
output N422; 
output N423; 
output N424; 
output N425; 
output N426; 
output N427; 
output N428; 
output N429; 
output N430; 
output N431; 
output N432; 
output N433; 
output N434; 
output N435; 
output N436; 
output N437; 
output N438; 
output N439; 
output N440; 
output N441; 
output N442; 
output N443; 
output N444; 
output N445; 
output N446; 
output N447; 
output N448; 
output N449; 
output N450; 
output N451; 
output N452; 
output N453; 
output N454; 
output N455; 
output N456; 
output N457; 
output N458; 
output N459; 
output N460; 
output N461; 
output N462; 
output N463; 
output N464; 
output N465; 
output N466; 
output N467; 
output N468; 
output N469; 
output N470; 
output N471; 
output N472; 
output N473; 
output N474; 
output N475; 
output N476; 
output N477; 

wire N7; 
wire N8; 
wire N9; 
wire N10; 
wire N11; 
wire N12; 
wire N13; 
wire N14; 
wire N15; 
wire N16; 
wire N17; 
wire N18; 
wire N19; 
wire N20; 
wire N21; 
wire N22; 
wire N23; 
wire N24; 
wire N25; 
wire N26; 
wire N27; 
wire N28; 
wire N29; 
wire N30; 
wire N31; 
wire N32; 
wire N33; 
wire N34; 
wire N35; 
wire N36; 
wire N37; 
wire N38; 
wire N39; 
wire N40; 
wire N41; 
wire N42; 
wire N43; 
wire N44; 
wire N45; 
wire N46; 
wire N47; 
wire N48; 
wire N49; 
wire N50; 
wire N51; 
wire N52; 
wire N53; 
wire N54; 
wire N55; 
wire N56; 
wire N57; 
wire N58; 
wire N59; 
wire N60; 
wire N61; 
wire N62; 
wire N63; 
wire N64; 
wire N65; 
wire N66; 
wire N67; 
wire N68; 
wire N69; 
wire N70; 
wire N71; 
wire N72; 
wire N73; 
wire N74; 
wire N75; 
wire N76; 
wire N77; 
wire N78; 
wire N79; 
wire N80; 
wire N81; 
wire N82; 
wire N83; 
wire N84; 
wire N85; 
wire N86; 
wire N87; 
wire N88; 
wire N89; 
wire N90; 
wire N91; 
wire N92; 
wire N93; 
wire N94; 
wire N95; 
wire N96; 
wire N97; 
wire N98; 
wire N99; 
wire N100; 
wire N101; 
wire N102; 
wire N103; 
wire N104; 
wire N105; 
wire N106; 
wire N107; 
wire N108; 
wire N109; 
wire N110; 
wire N111; 
wire N112; 
wire N113; 
wire N114; 
wire N115; 
wire N116; 
wire N117; 
wire N118; 
wire N119; 
wire N120; 
wire N121; 
wire N122; 
wire N123; 
wire N124; 
wire N125; 
wire N126; 
wire N127; 
wire N128; 
wire N129; 
wire N130; 
wire N131; 
wire N132; 
wire N133; 
wire N134; 
wire N135; 
wire N136; 
wire N137; 
wire N138; 
wire N139; 
wire N140; 
wire N141; 
wire N142; 
wire N143; 
wire N144; 
wire N145; 
wire N146; 
wire N147; 
wire N148; 
wire N149; 
wire N150; 
wire N151; 
wire N152; 
wire N153; 
wire N154; 
wire N155; 
wire N156; 
wire N157; 
wire N158; 
wire N159; 
wire N160; 
wire N161; 
wire N162; 
wire N163; 
wire N164; 
wire N165; 
wire N166; 
wire N167; 
wire N168; 
wire N169; 
wire N170; 
wire N171; 
wire N172; 
wire N173; 
wire N174; 
wire N175; 
wire N176; 
wire N177; 
wire N178; 
wire N179; 
wire N180; 
wire N181; 
wire N182; 
wire N183; 
wire N184; 
wire N185; 
wire N186; 
wire N187; 
wire N188; 
wire N189; 
wire N190; 
wire N191; 
wire N192; 
wire N193; 
wire N194; 
wire N195; 
wire N196; 
wire N197; 
wire N198; 
wire N199; 
wire N200; 
wire N201; 
wire N202; 
wire N203; 
wire N204; 
wire N205; 
wire N206; 
wire N207; 
wire N208; 
wire N209; 
wire N210; 
wire N211; 
wire N212; 
wire N213; 
wire N214; 
wire N215; 
wire N216; 
wire N217; 
wire N218; 
wire N219; 
wire N220; 
wire N221; 
wire N222; 
wire N223; 
wire N224; 
wire N225; 
wire N226; 
wire N227; 
wire N228; 
wire N229; 
wire N230; 
wire N231; 
wire N232; 
wire N233; 
wire N234; 
wire N235; 
wire N236; 
wire N237; 
wire N238; 
wire N239; 
wire N240; 
wire N241; 
wire N242; 
wire N243; 
wire N244; 
wire N245; 
wire N246; 
wire N247; 
wire N248; 
wire N249; 
wire N250; 
wire N251; 
wire N252; 
wire N253; 
wire N254; 
wire N255; 
wire N256; 
wire N257; 
wire N258; 
wire N259; 
wire N260; 
wire N261; 
wire N262; 
wire N263; 
wire N264; 
wire N265; 
wire N266; 
wire N267; 
wire N268; 
wire N269; 
wire N270; 
wire N271; 
wire N272; 
wire N273; 
wire N274; 
wire N275; 
wire N276; 
wire N277; 
wire N278; 
wire N279; 
wire N280; 
wire N281; 
wire N282; 
wire N283; 
wire N284; 
wire N285; 
wire N286; 
wire N287; 
wire N288; 
wire N289; 
wire N290; 
wire N291; 
wire N292; 
wire N293; 
wire N294; 
wire N295; 
wire N296; 
wire N297; 
wire N298; 
wire N299; 
wire N300; 
wire N301; 
wire N302; 
wire N303; 
wire N304; 
wire N305; 
wire N306; 
wire N307; 
wire N308; 
wire N309; 
wire N310; 
wire N311; 
wire N312; 
wire N313; 
wire N314; 
wire N315; 
wire N316; 
wire N317; 
wire N318; 
wire N319; 
wire N320; 
wire N321; 
wire N322; 
wire N323; 
wire N324; 
wire N325; 
wire N326; 
wire N327; 
wire N328; 
wire N329; 
wire N330; 
wire N331; 
wire N332; 
wire N333; 
wire N334; 
wire N335; 
wire N336; 
wire N337; 
wire N338; 
wire N339; 
wire N340; 
wire N341; 
wire N342; 
wire N343; 
wire N344; 
wire N345; 
wire N346; 
wire N347; 
wire N348; 
wire N349; 
wire N350; 
wire N351; 
wire N352; 
wire N353; 
wire N354; 
wire N355; 
wire N356; 
wire N357; 
wire N358; 
wire N359; 
wire N360; 
wire N361; 
wire N362; 
wire N363; 
wire N364; 
wire N365; 
wire N366; 
wire N367; 
wire N368; 
wire N369; 
wire N370; 
wire N371; 
wire N372; 
wire N373; 
wire N374; 
wire N375; 
wire N376; 
wire N377; 
wire N378; 
wire N379; 
wire N380; 
wire N381; 
wire N382; 
wire N383; 
wire N384; 
wire N385; 
wire N386; 
wire N387; 
wire N388; 
wire N389; 
wire N390; 
wire N391; 
wire N392; 
wire N393; 
wire N394; 
wire N395; 
wire N396; 
wire N397; 
wire N398; 
wire N399; 
wire N400; 
wire N401; 
wire N402; 
wire N403; 
wire N404; 
wire N405; 
wire N406; 
wire N407; 
wire N408; 
wire N409; 
wire N410; 
wire N411; 
wire N412; 
wire N413; 
wire N414; 

assign N7 = ~(N6); 
assign N8 = ~(N2); 
assign N9 = ~(N3); 
assign N10 = ~(N5); 
assign N11 = ~(N6); 
assign N12 = ~(N3); 
assign N13 = ~(N6); 
assign N14 = ~(N2); 
assign N15 = ~(N4); 
assign N16 = ~(N2); 
assign N17 = ~(N1); 
assign N18 = ~(N3); 
assign N19 = ~(N4); 
assign N20 = ~(N1); 
assign N21 = ~(N3); 
assign N22 = ~(N2); 
assign N23 = ~(N6); 
assign N24 = N18 & N4; 
assign N25 = ~(N16); 
assign N26 = ~(N2); 
assign N27 = ~(N4); 
assign N28 = ~(N8); 
assign N29 = ~(N17); 
assign N30 = ~(N4); 
assign N31 = N5 & N15; 
assign N32 = ~(N1); 
assign N33 = ~(N9); 
assign N34 = ~(N1); 
assign N35 = N7 & N12; 
assign N36 = N23 & N5; 
assign N37 = ~(N32); 
assign N38 = ~(N8); 
assign N39 = ~(N32); 
assign N40 = ~(N30); 
assign N41 = N15 & N33; 
assign N42 = N27 | N3; 
assign N43 = ~(N5); 
assign N44 = ~(N7); 
assign N45 = ~(N24); 
assign N46 = ~(N14); 
assign N47 = ~(N5); 
assign N48 = ~(N32); 
assign N49 = N28 & N33; 
assign N50 = ~(N30); 
assign N51 = N20 & N25; 
assign N52 = ~(N34); 
assign N53 = ~(N29); 
assign N54 = ~(N16); 
assign N55 = ~(N19); 
assign N56 = ~(N28); 
assign N57 = N11 & N26; 
assign N58 = ~(N9); 
assign N59 = ~(N10); 
assign N60 = ~(N21); 
assign N61 = ~(N12); 
assign N62 = ~(N31); 
assign N63 = ~(N18); 
assign N64 = N22 & N32; 
assign N65 = ~(N15); 
assign N66 = ~(N21); 
assign N67 = ~(N28); 
assign N68 = ~(N15); 
assign N69 = ~(N32); 
assign N70 = ~(N28); 
assign N71 = ~(N3); 
assign N72 = ~(N64); 
assign N73 = ~(N31); 
assign N74 = ~(N28); 
assign N75 = ~(N29); 
assign N76 = ~(N14); 
assign N77 = ~(N16); 
assign N78 = ~(N1); 
assign N79 = ~(N7); 
assign N80 = ~(N55); 
assign N81 = ~(N34); 
assign N82 = ~(N17); 
assign N83 = ~(N19); 
assign N84 = ~(N21); 
assign N85 = ~(N67); 
assign N86 = ~(N29); 
assign N87 = ~(N55); 
assign N88 = ~(N27); 
assign N89 = ~(N41); 
assign N90 = ~(N61); 
assign N91 = ~(N61); 
assign N92 = ~(N35); 
assign N93 = ~(N5); 
assign N94 = ~(N41); 
assign N95 = ~(N30); 
assign N96 = ~(N45); 
assign N97 = ~(N9); 
assign N98 = ~(N34); 
assign N99 = ~(N54); 
assign N100 = ~(N8); 
assign N101 = ~(N23); 
assign N102 = N9 | N29; 
assign N103 = ~(N25); 
assign N104 = ~(N42); 
assign N105 = ~(N26); 
assign N106 = ~(N6); 
assign N107 = ~(N33); 
assign N108 = ~(N64); 
assign N109 = ~(N19); 
assign N110 = ~(N33); 
assign N111 = ~(N24); 
assign N112 = ~(N17); 
assign N113 = ~(N48); 
assign N114 = ~(N31); 
assign N115 = ~(N22); 
assign N116 = ~(N11); 
assign N117 = ~(N35); 
assign N118 = ~(N37); 
assign N119 = ~(N38); 
assign N120 = N6 & N33; 
assign N121 = ~(N14); 
assign N122 = ~(N57); 
assign N123 = ~(N59); 
assign N124 = ~(N35); 
assign N125 = ~(N45); 
assign N126 = ~(N34); 
assign N127 = ~(N24); 
assign N128 = ~(N31); 
assign N129 = N24 | N18; 
assign N130 = ~(N26); 
assign N131 = ~(N12); 
assign N132 = ~(N9); 
assign N133 = ~(N18); 
assign N134 = ~(N46); 
assign N135 = ~(N35); 
assign N136 = ~(N11); 
assign N137 = ~(N68); 
assign N138 = ~(N37); 
assign N139 = ~(N64); 
assign N140 = ~(N51); 
assign N141 = ~(N49); 
assign N142 = ~(N28); 
assign N143 = ~(N69); 
assign N144 = ~(N35); 
assign N145 = ~(N31); 
assign N146 = ~(N7); 
assign N147 = ~(N25); 
assign N148 = ~(N52); 
assign N149 = ~(N47); 
assign N150 = ~(N9); 
assign N151 = ~(N12); 
assign N152 = ~(N14); 
assign N153 = ~(N50); 
assign N154 = ~(N22); 
assign N155 = ~(N20); 
assign N156 = ~(N27); 
assign N157 = ~(N20); 
assign N158 = ~(N62); 
assign N159 = ~(N37); 
assign N160 = ~(N46); 
assign N161 = ~(N36); 
assign N162 = ~(N52); 
assign N163 = ~(N11); 
assign N164 = ~(N23); 
assign N165 = ~(N38); 
assign N166 = ~(N24); 
assign N167 = ~(N51); 
assign N168 = ~(N63); 
assign N169 = ~(N62); 
assign N170 = ~(N40); 
assign N171 = ~(N17); 
assign N172 = ~(N48); 
assign N173 = ~(N63); 
assign N174 = ~(N46); 
assign N175 = ~(N42); 
assign N176 = ~(N37); 
assign N177 = ~(N10); 
assign N178 = ~(N30); 
assign N179 = ~(N46); 
assign N180 = ~(N55); 
assign N181 = ~(N65); 
assign N182 = ~(N62); 
assign N183 = ~(N12); 
assign N184 = ~(N59); 
assign N185 = ~(N64); 
assign N186 = ~(N46); 
assign N187 = ~(N29); 
assign N188 = ~(N17); 
assign N189 = ~(N22); 
assign N190 = ~(N45); 
assign N191 = ~(N53); 
assign N192 = ~(N50); 
assign N193 = ~(N8); 
assign N194 = ~(N13); 
assign N195 = ~(N58); 
assign N196 = ~(N39); 
assign N197 = ~(N63); 
assign N198 = ~(N57); 
assign N199 = ~(N24); 
assign N200 = ~(N47); 
assign N201 = ~(N21); 
assign N202 = N13 & N68; 
assign N203 = N21 | N46; 
assign N204 = ~(N8); 
assign N205 = ~(N66); 
assign N206 = ~(N53); 
assign N207 = ~(N36); 
assign N208 = ~(N66); 
assign N209 = ~(N67); 
assign N210 = ~(N37); 
assign N211 = ~(N26); 
assign N212 = ~(N62); 
assign N213 = ~(N56); 
assign N214 = ~(N47); 
assign N215 = ~(N26); 
assign N216 = ~(N67); 
assign N217 = ~(N11); 
assign N218 = ~(N54); 
assign N219 = ~(N34); 
assign N220 = ~(N16); 
assign N221 = ~(N40); 
assign N222 = ~(N39); 
assign N223 = ~(N44); 
assign N224 = ~(N44); 
assign N225 = ~(N134); 
assign N226 = N123 | N151; 
assign N227 = ~(N10); 
assign N228 = ~(N171); 
assign N229 = N87 | N158 | N159 | N212 | N23; 
assign N230 = N107 | N124 | N173; 
assign N231 = ~(N213); 
assign N232 = ~(N145); 
assign N233 = ~(N49); 
assign N234 = N113 & N205 & N221 & N201; 
assign N235 = ~(N53); 
assign N236 = N2 & N66; 
assign N237 = N82 & N137; 
assign N238 = N103 & N174 & N218; 
assign N239 = ~(N79); 
assign N240 = ~(N19); 
assign N241 = N89 & N156; 
assign N242 = N30 & N121 & N154 & N182 & N16; 
assign N243 = N14 | N44 | N59; 
assign N244 = N17 | N77 | N198 | N214; 
assign N245 = N93 | N241; 
assign N246 = ~(N53); 
assign N247 = ~(N41); 
assign N248 = ~(N52); 
assign N249 = N55 | N106 | N232 | N13; 
assign N250 = N165 & N201 & N72; 
assign N251 = ~(N65); 
assign N252 = N146 | N68; 
assign N253 = ~(N155); 
assign N254 = ~(N233); 
assign N255 = ~(N60); 
assign N256 = N127 & N15; 
assign N257 = ~(N52); 
assign N258 = ~(N16); 
assign N259 = N83 & N114 & N21; 
assign N260 = N197 | N236; 
assign N261 = ~(N232); 
assign N262 = ~(N50); 
assign N263 = N38 & N98 & N186; 
assign N264 = N133 & N55; 
assign N265 = N144 & N23; 
assign N266 = N4 & N235 & N43; 
assign N267 = ~(N211); 
assign N268 = N35 & N56; 
assign N269 = ~(N72); 
assign N270 = N189 & N25; 
assign N271 = N56 | N230; 
assign N272 = ~(N225); 
assign N273 = ~(N55); 
assign N274 = N220 | N23; 
assign N275 = N67 | N93; 
assign N276 = N32 | N7; 
assign N277 = ~(N40); 
assign N278 = N51 & N50; 
assign N279 = ~(N232); 
assign N280 = ~(N146); 
assign N281 = ~(N105); 
assign N282 = N188 | N195; 
assign N283 = ~(N96); 
assign N284 = ~(N233); 
assign N285 = ~(N51); 
assign N286 = ~(N27); 
assign N287 = ~(N15); 
assign N288 = N53 | N68 | N63; 
assign N289 = ~(N74); 
assign N290 = ~(N175); 
assign N291 = N29 | N108 | N244; 
assign N292 = ~(N22); 
assign N293 = ~(N121); 
assign N294 = ~(N1); 
assign N295 = ~(N243); 
assign N296 = ~(N13); 
assign N297 = N33 | N84 | N118 | N210 | N288 | N116; 
assign N298 = N25 & N78 & N90 & N204 & N228 & N238 & N261 & N292; 
assign N299 = N34 & N58 & N85 & N97 & N132 & N162 & N194 & N209; 
assign N300 = N26 | N91 | N153 | N164 | N177 | N225 | N246 | N267; 
assign N301 = N31 | N37 | N40 | N139 | N148 | N161 | N187 | N277; 
assign N302 = N12 & N81 & N112 & N136 & N196 & N207 & N251 & N270; 
assign N303 = N19 | N80 | N101 | N168 | N248 | N27; 
assign N304 = ~(N64); 
assign N305 = ~(N125); 
assign N306 = N71 | N135; 
assign N307 = N170 | N224; 
assign N308 = N104 | N183 | N191 | N219 | N50; 
assign N309 = ~(N264); 
assign N310 = N36 | N140 | N230; 
assign N311 = N92 | N237 | N231; 
assign N312 = ~(N276); 
assign N313 = ~(N120); 
assign N314 = N59 & N147 & N176 & N214; 
assign N315 = N141 & N157 & N233; 
assign N316 = N275 & N175; 
assign N317 = ~(N83); 
assign N318 = ~(N268); 
assign N319 = ~(N54); 
assign N320 = N61 & N88 & N211 & N213; 
assign N321 = N52 & N86 & N131 & N245; 
assign N322 = N43 | N301; 
assign N323 = N60 | N243 | N69; 
assign N324 = N240 | N62; 
assign N325 = ~(N59); 
assign N326 = N102 | N203 | N173; 
assign N327 = N122 | N128 | N252 | N293; 
assign N328 = N119 | N217 | N262 | N240 | N287; 
assign N329 = N129 & N152 & N272 & N127; 
assign N330 = N50 | N63 | N109 | N179 | N215 | N241; 
assign N331 = N70 | N200 | N208 | N306 | N20; 
assign N332 = N130 & N190 & N227 & N229; 
assign N333 = N45 | N75 | N202 | N250 | N313 | N178; 
assign N334 = N47 & N111 & N273 & N20 & N314; 
assign N335 = N41 | N42 | N48 | N94 | N160 | N40; 
assign N336 = N39 & N62 & N69 & N73 & N95 & N138 & N167 & N309; 
assign N337 = N99 | N169 | N242 | N281; 
assign N338 = ~(N298); 
assign N339 = N65 | N178 | N216 | N236 | N285; 
assign N340 = N110 | N195 | N320; 
assign N341 = N256 & N286 & N291 & N323 & N65; 
assign N342 = N192 & N223 & N254 & N299 & N30; 
assign N343 = N172 & N224; 
assign N344 = N116 & N135 & N185 & N231 & N269 & N80; 
assign N345 = N304 & N278; 
assign N346 = ~(N180); 
assign N347 = N100 & N166 & N199 & N222 & N41; 
assign N348 = N266 | N326 | N18; 
assign N349 = N171 & N184 & N183 & N328; 
assign N350 = N115 & N175 & N181; 
assign N351 = N126 & N193 & N27; 
assign N352 = N206 | N241 | N315; 
assign N353 = N302 | N83; 
assign N354 = N303 & N165; 
assign N355 = N253 | N259 | N271 | N20; 
assign N356 = N308 & N321 & N239; 
assign N357 = ~(N164); 
assign N358 = N76 | N143 | N249 | N289 | N297 | N40; 
assign N359 = N117 | N239 | N44; 
assign N360 = N105 | N142 | N149 | N150 | N163 | N233 | N263 | N265; 
assign N361 = N229 & N244; 
assign N362 = N226 | N290 | N294; 
assign N363 = ~(N113); 
assign N364 = N344 & N61; 
assign N365 = N356 | N104; 
assign N366 = ~(N226); 
assign N367 = ~(N274); 
assign N368 = ~(N196); 
assign N369 = ~(N255); 
assign N370 = ~(N122); 
assign N371 = ~(N352); 
assign N372 = N260 | N108; 
assign N373 = N317 | N318 | N229; 
assign N374 = N234 | N336 | N51; 
assign N375 = N305 | N237 | N282; 
assign N376 = N257 & N78; 
assign N377 = ~(N346); 
assign N378 = N350 | N374 | N241; 
assign N379 = N280 & N362 & N371; 
assign N380 = N316 | N330 | N345 | N353 | N367 | N235; 
assign N381 = N331 & N14; 
assign N382 = N373 | N232; 
assign N383 = N284 | N346; 
assign N384 = N247 & N279 & N298 & N351 & N354; 
assign N385 = N300 | N327 | N18; 
assign N386 = N283 & N339 & N349; 
assign N387 = N381 | N44; 
assign N388 = ~(N244); 
assign N389 = ~(N227); 
assign N390 = N359 & N196; 
assign N391 = N357 & N363 & N382 & N386; 
assign N392 = N324 | N369; 
assign N393 = ~(N236); 
assign N394 = N343 & N230; 
assign N395 = N370 & N38; 
assign N396 = ~(N8); 
assign N397 = ~(N141); 
assign N398 = ~(N176); 
assign N399 = ~(N361); 
assign N400 = N341 | N360; 
assign N401 = ~(N382); 
assign N402 = ~(N305); 
assign N403 = ~(N68); 
assign N404 = ~(N385); 
assign N405 = N319 & N25; 
assign N406 = ~(N217); 
assign N407 = N375 | N239; 
assign N408 = ~(N57); 
assign N409 = N338 | N347 | N378 | N213; 
assign N410 = ~(N83); 
assign N411 = ~(N66); 
assign N412 = ~(N13); 
assign N413 = ~(N277); 
assign N414 = N335 & N376 & N47; 
assign N415 = N333 | N368 | N402; 
assign N416 = ~(N351); 
assign N417 = ~(N393); 
assign N418 = N332 | N348; 
assign N419 = ~(N334); 
assign N420 = N372 | N410; 
assign N421 = ~(N345); 
assign N422 = N388 | N397 | N401; 
assign N423 = ~(N405); 
assign N424 = N379 | N399; 
assign N425 = ~(N319); 
assign N426 = ~(N282); 
assign N427 = ~(N412); 
assign N428 = ~(N329); 
assign N429 = N390 & N408; 
assign N430 = N377 & N414; 
assign N431 = ~(N342); 
assign N432 = N392 | N400; 
assign N433 = ~(N282); 
assign N434 = ~(N53); 
assign N435 = ~(N295); 
assign N436 = ~(N300); 
assign N437 = ~(N342); 
assign N438 = ~(N409); 
assign N439 = ~(N11); 
assign N440 = ~(N364); 
assign N441 = N322 | N310; 
assign N442 = ~(N411); 
assign N443 = ~(N217); 
assign N444 = ~(N347); 
assign N445 = N389 & N396 & N296; 
assign N446 = ~(N299); 
assign N447 = ~(N332); 
assign N448 = ~(N355); 
assign N449 = ~(N151); 
assign N450 = N312 & N393; 
assign N451 = ~(N307); 
assign N452 = ~(N52); 
assign N453 = N365 & N380; 
assign N454 = ~(N394); 
assign N455 = ~(N384); 
assign N456 = ~(N328); 
assign N457 = ~(N231); 
assign N458 = ~(N395); 
assign N459 = ~(N233); 
assign N460 = ~(N350); 
assign N461 = ~(N22); 
assign N462 = ~(N414); 
assign N463 = N383 & N407; 
assign N464 = ~(N346); 
assign N465 = ~(N340); 
assign N466 = N340 | N406; 
assign N467 = N361 & N387; 
assign N468 = N337 | N358 | N404; 
assign N469 = ~(N395); 
assign N470 = ~(N239); 
assign N471 = ~(N63); 
assign N472 = ~(N413); 
assign N473 = ~(N258); 
assign N474 = N385 | N391 | N398; 
assign N475 = ~(N222); 
assign N476 = N325 | N366; 
assign N477 = N311 | N403; 
endmodule
