module Depth_10_20_Nodes_200_400_S005 (N1, N2, N3, N4, N5, N6, N7, N8, N9, N306, N307, N308, N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319, N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330, N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341, N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352, N353, N354);

input N1; 
input N2; 
input N3; 
input N4; 
input N5; 
input N6; 
input N7; 
input N8; 
input N9; 

output N306; 
output N307; 
output N308; 
output N309; 
output N310; 
output N311; 
output N312; 
output N313; 
output N314; 
output N315; 
output N316; 
output N317; 
output N318; 
output N319; 
output N320; 
output N321; 
output N322; 
output N323; 
output N324; 
output N325; 
output N326; 
output N327; 
output N328; 
output N329; 
output N330; 
output N331; 
output N332; 
output N333; 
output N334; 
output N335; 
output N336; 
output N337; 
output N338; 
output N339; 
output N340; 
output N341; 
output N342; 
output N343; 
output N344; 
output N345; 
output N346; 
output N347; 
output N348; 
output N349; 
output N350; 
output N351; 
output N352; 
output N353; 
output N354; 

wire N10; 
wire N11; 
wire N12; 
wire N13; 
wire N14; 
wire N15; 
wire N16; 
wire N17; 
wire N18; 
wire N19; 
wire N20; 
wire N21; 
wire N22; 
wire N23; 
wire N24; 
wire N25; 
wire N26; 
wire N27; 
wire N28; 
wire N29; 
wire N30; 
wire N31; 
wire N32; 
wire N33; 
wire N34; 
wire N35; 
wire N36; 
wire N37; 
wire N38; 
wire N39; 
wire N40; 
wire N41; 
wire N42; 
wire N43; 
wire N44; 
wire N45; 
wire N46; 
wire N47; 
wire N48; 
wire N49; 
wire N50; 
wire N51; 
wire N52; 
wire N53; 
wire N54; 
wire N55; 
wire N56; 
wire N57; 
wire N58; 
wire N59; 
wire N60; 
wire N61; 
wire N62; 
wire N63; 
wire N64; 
wire N65; 
wire N66; 
wire N67; 
wire N68; 
wire N69; 
wire N70; 
wire N71; 
wire N72; 
wire N73; 
wire N74; 
wire N75; 
wire N76; 
wire N77; 
wire N78; 
wire N79; 
wire N80; 
wire N81; 
wire N82; 
wire N83; 
wire N84; 
wire N85; 
wire N86; 
wire N87; 
wire N88; 
wire N89; 
wire N90; 
wire N91; 
wire N92; 
wire N93; 
wire N94; 
wire N95; 
wire N96; 
wire N97; 
wire N98; 
wire N99; 
wire N100; 
wire N101; 
wire N102; 
wire N103; 
wire N104; 
wire N105; 
wire N106; 
wire N107; 
wire N108; 
wire N109; 
wire N110; 
wire N111; 
wire N112; 
wire N113; 
wire N114; 
wire N115; 
wire N116; 
wire N117; 
wire N118; 
wire N119; 
wire N120; 
wire N121; 
wire N122; 
wire N123; 
wire N124; 
wire N125; 
wire N126; 
wire N127; 
wire N128; 
wire N129; 
wire N130; 
wire N131; 
wire N132; 
wire N133; 
wire N134; 
wire N135; 
wire N136; 
wire N137; 
wire N138; 
wire N139; 
wire N140; 
wire N141; 
wire N142; 
wire N143; 
wire N144; 
wire N145; 
wire N146; 
wire N147; 
wire N148; 
wire N149; 
wire N150; 
wire N151; 
wire N152; 
wire N153; 
wire N154; 
wire N155; 
wire N156; 
wire N157; 
wire N158; 
wire N159; 
wire N160; 
wire N161; 
wire N162; 
wire N163; 
wire N164; 
wire N165; 
wire N166; 
wire N167; 
wire N168; 
wire N169; 
wire N170; 
wire N171; 
wire N172; 
wire N173; 
wire N174; 
wire N175; 
wire N176; 
wire N177; 
wire N178; 
wire N179; 
wire N180; 
wire N181; 
wire N182; 
wire N183; 
wire N184; 
wire N185; 
wire N186; 
wire N187; 
wire N188; 
wire N189; 
wire N190; 
wire N191; 
wire N192; 
wire N193; 
wire N194; 
wire N195; 
wire N196; 
wire N197; 
wire N198; 
wire N199; 
wire N200; 
wire N201; 
wire N202; 
wire N203; 
wire N204; 
wire N205; 
wire N206; 
wire N207; 
wire N208; 
wire N209; 
wire N210; 
wire N211; 
wire N212; 
wire N213; 
wire N214; 
wire N215; 
wire N216; 
wire N217; 
wire N218; 
wire N219; 
wire N220; 
wire N221; 
wire N222; 
wire N223; 
wire N224; 
wire N225; 
wire N226; 
wire N227; 
wire N228; 
wire N229; 
wire N230; 
wire N231; 
wire N232; 
wire N233; 
wire N234; 
wire N235; 
wire N236; 
wire N237; 
wire N238; 
wire N239; 
wire N240; 
wire N241; 
wire N242; 
wire N243; 
wire N244; 
wire N245; 
wire N246; 
wire N247; 
wire N248; 
wire N249; 
wire N250; 
wire N251; 
wire N252; 
wire N253; 
wire N254; 
wire N255; 
wire N256; 
wire N257; 
wire N258; 
wire N259; 
wire N260; 
wire N261; 
wire N262; 
wire N263; 
wire N264; 
wire N265; 
wire N266; 
wire N267; 
wire N268; 
wire N269; 
wire N270; 
wire N271; 
wire N272; 
wire N273; 
wire N274; 
wire N275; 
wire N276; 
wire N277; 
wire N278; 
wire N279; 
wire N280; 
wire N281; 
wire N282; 
wire N283; 
wire N284; 
wire N285; 
wire N286; 
wire N287; 
wire N288; 
wire N289; 
wire N290; 
wire N291; 
wire N292; 
wire N293; 
wire N294; 
wire N295; 
wire N296; 
wire N297; 
wire N298; 
wire N299; 
wire N300; 
wire N301; 
wire N302; 
wire N303; 
wire N304; 
wire N305; 

assign N10 = ~(N4); 
assign N11 = ~(N4); 
assign N12 = ~(N2); 
assign N13 = ~(N8); 
assign N14 = N4 & N5; 
assign N15 = ~(N11); 
assign N16 = ~(N8); 
assign N17 = N9 | N10; 
assign N18 = ~(N4); 
assign N19 = ~(N6); 
assign N20 = ~(N4); 
assign N21 = ~(N10); 
assign N22 = ~(N10); 
assign N23 = ~(N10); 
assign N24 = ~(N12); 
assign N25 = ~(N5); 
assign N26 = ~(N2); 
assign N27 = ~(N13); 
assign N28 = ~(N13); 
assign N29 = ~(N12); 
assign N30 = ~(N3); 
assign N31 = ~(N11); 
assign N32 = ~(N5); 
assign N33 = ~(N1); 
assign N34 = ~(N13); 
assign N35 = ~(N13); 
assign N36 = ~(N6); 
assign N37 = ~(N14); 
assign N38 = ~(N12); 
assign N39 = ~(N11); 
assign N40 = ~(N4); 
assign N41 = ~(N5); 
assign N42 = ~(N25); 
assign N43 = ~(N2); 
assign N44 = ~(N23); 
assign N45 = ~(N5); 
assign N46 = ~(N11); 
assign N47 = ~(N30); 
assign N48 = N33 & N3; 
assign N49 = ~(N13); 
assign N50 = ~(N9); 
assign N51 = ~(N6); 
assign N52 = ~(N24); 
assign N53 = ~(N6); 
assign N54 = N36 & N17; 
assign N55 = ~(N9); 
assign N56 = ~(N19); 
assign N57 = N15 | N9; 
assign N58 = ~(N12); 
assign N59 = ~(N30); 
assign N60 = ~(N3); 
assign N61 = ~(N20); 
assign N62 = ~(N20); 
assign N63 = ~(N36); 
assign N64 = ~(N10); 
assign N65 = ~(N56); 
assign N66 = ~(N3); 
assign N67 = N5 | N26; 
assign N68 = N29 | N63 | N9; 
assign N69 = ~(N12); 
assign N70 = N57 & N41; 
assign N71 = N46 | N56; 
assign N72 = N2 | N13; 
assign N73 = N50 & N44; 
assign N74 = ~(N26); 
assign N75 = N61 & N8; 
assign N76 = ~(N14); 
assign N77 = ~(N20); 
assign N78 = ~(N67); 
assign N79 = ~(N73); 
assign N80 = ~(N14); 
assign N81 = ~(N20); 
assign N82 = ~(N56); 
assign N83 = N71 & N8; 
assign N84 = ~(N71); 
assign N85 = ~(N74); 
assign N86 = N24 | N39; 
assign N87 = ~(N65); 
assign N88 = N52 & N66; 
assign N89 = N69 & N48; 
assign N90 = N62 | N34; 
assign N91 = ~(N11); 
assign N92 = ~(N33); 
assign N93 = ~(N41); 
assign N94 = ~(N24); 
assign N95 = N26 & N73; 
assign N96 = ~(N91); 
assign N97 = ~(N2); 
assign N98 = ~(N8); 
assign N99 = N81 & N83; 
assign N100 = N3 & N22 & N42 & N45 & N84 & N93; 
assign N101 = ~(N85); 
assign N102 = ~(N81); 
assign N103 = ~(N14); 
assign N104 = N19 & N18; 
assign N105 = ~(N54); 
assign N106 = ~(N41); 
assign N107 = N23 & N87 & N99; 
assign N108 = N98 | N20; 
assign N109 = N18 & N93; 
assign N110 = ~(N93); 
assign N111 = ~(N99); 
assign N112 = ~(N51); 
assign N113 = ~(N100); 
assign N114 = ~(N95); 
assign N115 = ~(N81); 
assign N116 = ~(N69); 
assign N117 = ~(N74); 
assign N118 = ~(N20); 
assign N119 = ~(N15); 
assign N120 = ~(N80); 
assign N121 = ~(N6); 
assign N122 = ~(N7); 
assign N123 = ~(N97); 
assign N124 = N44 & N68 & N76; 
assign N125 = ~(N23); 
assign N126 = ~(N93); 
assign N127 = ~(N67); 
assign N128 = N16 & N77 & N7; 
assign N129 = ~(N44); 
assign N130 = N8 & N27; 
assign N131 = N122 | N121; 
assign N132 = ~(N30); 
assign N133 = ~(N31); 
assign N134 = ~(N60); 
assign N135 = ~(N31); 
assign N136 = ~(N10); 
assign N137 = ~(N52); 
assign N138 = ~(N98); 
assign N139 = ~(N44); 
assign N140 = N12 & N106 & N9; 
assign N141 = ~(N123); 
assign N142 = ~(N116); 
assign N143 = N78 | N89 | N125 | N63; 
assign N144 = ~(N89); 
assign N145 = N40 & N59 & N111; 
assign N146 = ~(N132); 
assign N147 = N88 & N128 & N29; 
assign N148 = N37 & N50; 
assign N149 = N72 | N96; 
assign N150 = ~(N84); 
assign N151 = N14 & N58 & N115 & N99; 
assign N152 = N17 | N54 | N136; 
assign N153 = ~(N91); 
assign N154 = N66 | N91 | N129; 
assign N155 = ~(N140); 
assign N156 = N133 | N124; 
assign N157 = N129 & N130; 
assign N158 = N70 & N142 & N34; 
assign N159 = N1 & N75; 
assign N160 = N7 | N64 | N82 | N113 | N123 | N93; 
assign N161 = N105 & N149 & N150 & N17; 
assign N162 = N90 | N118 | N152; 
assign N163 = N103 | N100; 
assign N164 = ~(N6); 
assign N165 = ~(N133); 
assign N166 = ~(N98); 
assign N167 = ~(N96); 
assign N168 = ~(N63); 
assign N169 = N11 & N85; 
assign N170 = ~(N18); 
assign N171 = N114 | N154 | N96; 
assign N172 = ~(N53); 
assign N173 = N49 & N143 & N105; 
assign N174 = ~(N65); 
assign N175 = N76 | N52; 
assign N176 = ~(N97); 
assign N177 = ~(N35); 
assign N178 = ~(N36); 
assign N179 = ~(N7); 
assign N180 = ~(N100); 
assign N181 = ~(N100); 
assign N182 = ~(N41); 
assign N183 = N120 & N145; 
assign N184 = ~(N80); 
assign N185 = ~(N69); 
assign N186 = ~(N152); 
assign N187 = ~(N99); 
assign N188 = N101 | N96; 
assign N189 = ~(N133); 
assign N190 = ~(N80); 
assign N191 = ~(N29); 
assign N192 = N130 | N65; 
assign N193 = ~(N112); 
assign N194 = ~(N54); 
assign N195 = ~(N139); 
assign N196 = ~(N37); 
assign N197 = N28 | N116 | N96; 
assign N198 = N38 & N178 & N146; 
assign N199 = ~(N78); 
assign N200 = N41 | N47 | N144 | N172 | N176 | N56; 
assign N201 = N48 | N51; 
assign N202 = N25 | N32; 
assign N203 = N27 | N195 | N87; 
assign N204 = ~(N21); 
assign N205 = N34 & N85 & N98; 
assign N206 = N43 & N138 & N49; 
assign N207 = ~(N109); 
assign N208 = N97 | N206 | N68; 
assign N209 = N147 & N152; 
assign N210 = N67 & N163 & N203 & N73; 
assign N211 = ~(N45); 
assign N212 = N74 | N32; 
assign N213 = N55 & N188 & N1; 
assign N214 = ~(N71); 
assign N215 = N95 | N99 | N126 | N180 | N97; 
assign N216 = N75 | N92 | N135 | N189 | N1; 
assign N217 = ~(N194); 
assign N218 = N117 | N159; 
assign N219 = N79 | N124 | N161 | N196 | N143; 
assign N220 = ~(N155); 
assign N221 = ~(N151); 
assign N222 = N167 & N150; 
assign N223 = ~(N137); 
assign N224 = N164 | N175 | N136; 
assign N225 = N134 & N139 & N158 & N94; 
assign N226 = N187 & N207 & N44; 
assign N227 = N109 & N156; 
assign N228 = N80 & N157 & N152; 
assign N229 = N212 & N226 & N65; 
assign N230 = N104 & N124; 
assign N231 = N186 | N40; 
assign N232 = ~(N97); 
assign N233 = N211 | N66; 
assign N234 = ~(N206); 
assign N235 = ~(N213); 
assign N236 = ~(N48); 
assign N237 = ~(N131); 
assign N238 = ~(N225); 
assign N239 = ~(N139); 
assign N240 = N102 | N132 | N96; 
assign N241 = ~(N95); 
assign N242 = N110 | N111 | N121 | N127; 
assign N243 = N136 | N104; 
assign N244 = ~(N114); 
assign N245 = ~(N130); 
assign N246 = ~(N98); 
assign N247 = N94 | N117; 
assign N248 = N86 | N84; 
assign N249 = N199 | N143; 
assign N250 = ~(N95); 
assign N251 = ~(N43); 
assign N252 = ~(N132); 
assign N253 = ~(N137); 
assign N254 = ~(N111); 
assign N255 = N137 & N185 & N139; 
assign N256 = ~(N90); 
assign N257 = ~(N7); 
assign N258 = ~(N46); 
assign N259 = ~(N142); 
assign N260 = ~(N135); 
assign N261 = ~(N90); 
assign N262 = ~(N130); 
assign N263 = ~(N128); 
assign N264 = ~(N14); 
assign N265 = ~(N218); 
assign N266 = N201 | N109; 
assign N267 = N245 & N83; 
assign N268 = N230 | N239; 
assign N269 = N202 & N105; 
assign N270 = N140 & N150; 
assign N271 = ~(N22); 
assign N272 = N192 & N65; 
assign N273 = ~(N57); 
assign N274 = ~(N160); 
assign N275 = ~(N163); 
assign N276 = N198 | N228 | N133; 
assign N277 = N152 & N234 & N45; 
assign N278 = ~(N144); 
assign N279 = N220 | N86; 
assign N280 = ~(N85); 
assign N281 = N170 | N29; 
assign N282 = N227 | N244 | N148; 
assign N283 = ~(N161); 
assign N284 = N193 | N126; 
assign N285 = N145 | N261 | N113; 
assign N286 = N256 | N60; 
assign N287 = ~(N79); 
assign N288 = N217 & N221 & N223 & N107; 
assign N289 = N243 | N147; 
assign N290 = ~(N148); 
assign N291 = ~(N66); 
assign N292 = N253 | N1; 
assign N293 = ~(N58); 
assign N294 = ~(N107); 
assign N295 = N100 & N263 & N73; 
assign N296 = ~(N219); 
assign N297 = N131 | N174 | N17; 
assign N298 = N119 & N127 & N148 & N184 & N240 & N252 & N254 & N260; 
assign N299 = N200 & N205 & N222 & N233 & N255 & N265 & N272 & N283; 
assign N300 = N224 | N249 | N271 | N284 | N276 | N293; 
assign N301 = N204 | N237 | N241 | N290 | N294 | N109; 
assign N302 = N112 | N146 | N169 | N295; 
assign N303 = N183 | N246 | N248 | N275 | N278; 
assign N304 = N208 & N218 & N229 & N247 & N270 & N277 & N280 & N296 & N282; 
assign N305 = N108 | N173 | N177 | N262 | N264 | N274 | N143; 
assign N306 = ~(N19); 
assign N307 = N279 | N287; 
assign N308 = ~(N105); 
assign N309 = N171 & N266; 
assign N310 = ~(N209); 
assign N311 = ~(N218); 
assign N312 = N179 & N269; 
assign N313 = ~(N239); 
assign N314 = ~(N37); 
assign N315 = ~(N197); 
assign N316 = ~(N126); 
assign N317 = ~(N286); 
assign N318 = ~(N216); 
assign N319 = N162 | N210 | N238 | N257; 
assign N320 = N242 | N273; 
assign N321 = N235 & N259; 
assign N322 = ~(N232); 
assign N323 = ~(N281); 
assign N324 = ~(N302); 
assign N325 = ~(N190); 
assign N326 = ~(N247); 
assign N327 = ~(N156); 
assign N328 = N299 & N285 & N292; 
assign N329 = ~(N304); 
assign N330 = ~(N141); 
assign N331 = ~(N267); 
assign N332 = N191 | N250; 
assign N333 = N166 & N258; 
assign N334 = N168 | N215; 
assign N335 = N301 | N303; 
assign N336 = ~(N231); 
assign N337 = ~(N304); 
assign N338 = ~(N300); 
assign N339 = ~(N153); 
assign N340 = ~(N15); 
assign N341 = ~(N153); 
assign N342 = ~(N291); 
assign N343 = ~(N145); 
assign N344 = N297 & N298; 
assign N345 = ~(N214); 
assign N346 = ~(N95); 
assign N347 = N165 | N251; 
assign N348 = N182 & N288 & N305; 
assign N349 = ~(N289); 
assign N350 = N236 & N268; 
assign N351 = ~(N181); 
assign N352 = ~(N97); 
assign N353 = ~(N88); 
assign N354 = ~(N166); 
endmodule
